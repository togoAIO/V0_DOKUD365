[{"log_codes":["UidNotFound"],"type":"Conceptual","source_relative_path":"ProcessDoku/01_CoreProcesses/01_03_Sales/Customer.md","output":{".html":{"relative_path":"ProcessDoku/01_CoreProcesses/01_03_Sales/Customer.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\whgw2ehc.c4q","hash":"j37StSW9xyc1v54fgIUoeA=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"customer\" sourcefile=\"ProcessDoku/01_CoreProcesses/01_03_Sales/Customer.md\" sourcestartlinenumber=\"5\">Customer</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/01_CoreProcesses/01_03_Sales/Guideline.md","output":{".html":{"relative_path":"ProcessDoku/01_CoreProcesses/01_03_Sales/Guideline.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\lgn44wd4.p2w","hash":"/z3EufMOMNa0D1BOJxIxFQ=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"guideline\" sourcefile=\"ProcessDoku/01_CoreProcesses/01_03_Sales/Guideline.md\" sourcestartlinenumber=\"5\">Guideline</h1>"},{"log_codes":["InvalidFileLink"],"type":"Conceptual","source_relative_path":"ProcessDoku/01_CoreProcesses/01_03_Sales/Sales.md","output":{".html":{"relative_path":"ProcessDoku/01_CoreProcesses/01_03_Sales/Sales.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\4rebvovl.mfi","hash":"lIgwqXmsvQykFHuyt8VDsA=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"sales-overview\" sourcefile=\"ProcessDoku/01_CoreProcesses/01_03_Sales/Sales.md\" sourcestartlinenumber=\"1\">Sales overview</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/01_CoreProcesses/01_01_CRM/CRM.md","output":{".html":{"relative_path":"ProcessDoku/01_CoreProcesses/01_01_CRM/CRM.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\jghujqhm.ute","hash":"rBKpqLbiJpFqwEj/U2yDBw=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"crm\" sourcefile=\"ProcessDoku/01_CoreProcesses/01_01_CRM/CRM.md\" sourcestartlinenumber=\"1\">CRM</h1>"},{"log_codes":["InvalidFileLink"],"type":"Conceptual","source_relative_path":"ProcessDoku/01_CoreProcesses/CoreProcesses_Overview.md","output":{".html":{"relative_path":"ProcessDoku/01_CoreProcesses/CoreProcesses_Overview.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\lroje5el.skl","hash":"RS4wOdG5IQmShAnW0U0uUw=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"core-processes-overview\" sourcefile=\"ProcessDoku/01_CoreProcesses/CoreProcesses_Overview.md\" sourcestartlinenumber=\"1\">Core Processes Overview</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/create-legal-entity.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/create-legal-entity.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\1ztu3k1q.kgm","hash":"6vlyi0Xomt2on2S+xUmnbw=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"create-a-legal-entity\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/create-legal-entity.md\" sourcestartlinenumber=\"25\">Erstellen Sie eine juristische Person</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/configure-global-address-book.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/configure-global-address-book.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\2vwfcjma.5cd","hash":"WRtrHlSVy0hvAH0HnBrD3w=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"configure-the-global-address-book\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/configure-global-address-book.md\" sourcestartlinenumber=\"25\">Konfigurieren des globalen Adressbuchs</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/qa-address-books.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/qa-address-books.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\slrffhox.nei","hash":"W+jSIhCMnKCyXrifhVSh9A=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"address-books-faq\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/organization-administration/qa-address-books.md\" sourcestartlinenumber=\"27\">FAQs zu Adressbüchern</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/plan-organizational-hierarchy.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/plan-organizational-hierarchy.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\nweihroa.odv","hash":"uftKBFsX5dptsN2ovCeqXQ=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"plan-your-organizational-hierarchy\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/organization-administration/plan-organizational-hierarchy.md\" sourcestartlinenumber=\"27\">Planen Ihrer Organisationshierarchie</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/configure-parallel-branch-workflow.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/configure-parallel-branch-workflow.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\qjne5vub.ypp","hash":"PQAWEAvn05p5fvJ+eNNsew=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"configure-parallel-branches-in-a-workflow\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/organization-administration/configure-parallel-branch-workflow.md\" sourcestartlinenumber=\"26\">Konfigurieren paralleler Verzweigungen in einem Workflow</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/configure-parallel-activity-workflow.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/configure-parallel-activity-workflow.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\tsyfggdc.px1","hash":"JHevHOUkJIcbu74vLnojSg=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"configure-parallel-activities-in-a-workflow\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/organization-administration/configure-parallel-activity-workflow.md\" sourcestartlinenumber=\"26\">Konfigurieren paralleler Aktivitäten in einem Workflow</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/configure-manual-decision-workflow.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/configure-manual-decision-workflow.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\caskrz5k.zpv","hash":"jcHAONu7hthfjDACMl0r9w=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"configure-manual-decisions-in-a-workflow\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/organization-administration/configure-manual-decision-workflow.md\" sourcestartlinenumber=\"26\">Manuellen Entscheidungen in einem Workflow konfigurieren</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/configure-automated-task-workflow.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/configure-automated-task-workflow.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\mojbcdzi.kgx","hash":"NiTvi5CF6xA8kBV+PdTt2g=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"configure-automated-tasks-in-a-workflow\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/organization-administration/configure-automated-task-workflow.md\" sourcestartlinenumber=\"26\">Konfigurieren von automatisierten Aufgaben in einem Workflow</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/hr/tasks/hire-candidate-through-recruiting.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/hr/tasks/hire-candidate-through-recruiting.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\cpbywrgk.zk0","hash":"9Mp7C9kfP7ot8FAKAQI/TQ=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"hiring-candidate-through-recruiting\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/hr/tasks/hire-candidate-through-recruiting.md\" sourcestartlinenumber=\"25\">Kandidaten über Rekrutierung einstellen</h1>"},{"log_codes":["InvalidFileLink"],"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/hr/hr-landing-page.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/hr/hr-landing-page.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\3xgvkwkd.wmx","hash":"s/KtYizr2D6GA4r1bvPqVA=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"human-resources-overview\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/hr/hr-landing-page.md\" sourcestartlinenumber=\"25\">Personalwesen – Übersicht</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/user-defined-fields.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/user-defined-fields.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\vozctahw.2rc","hash":"z9AqZsHQ536O3q4j2ksu6w=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"create-and-work-with-custom-fields\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/get-started/user-defined-fields.md\" sourcestartlinenumber=\"25\">Erstellen von und Arbeiten mit benutzerdefinierten Feldern</h1>"},{"log_codes":["InvalidFileLink"],"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/personalize-user-experience.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/personalize-user-experience.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\t3h1r1yy.dkr","hash":"54eeJPD1DnkZ8hh3yKldcw=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"personalize-the-user-experience\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/get-started/personalize-user-experience.md\" sourcestartlinenumber=\"27\">Die Benutzerumgebung personalisieren</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/feature-management/feature-management-overview.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/feature-management/feature-management-overview.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\4gce4f4w.f0n","hash":"empAlTFI5tC4xBNd+lh7xg=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"feature-management-overview\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/get-started/feature-management/feature-management-overview.md\" sourcestartlinenumber=\"27\">Funktionsverwaltung – Übersicht</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/use-lookups-to-find-information.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/use-lookups-to-find-information.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\ygmmaoey.vym","hash":"7CgFQN/EIvb3TRvVrMFwew=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"find-information-by-using-lookups\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/get-started/use-lookups-to-find-information.md\" sourcestartlinenumber=\"26\">Informationen per Suchen finden</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/configure-filter-workspaces.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/configure-filter-workspaces.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\eyjy20qm.m4p","hash":"kiqGCrFtPmTAr2brxM0bbA=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"configure-and-filter-workspaces\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/get-started/configure-filter-workspaces.md\" sourcestartlinenumber=\"27\">Arbeitsbereiche konfigurieren und Filtern</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/alert-email-notifications.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/alert-email-notifications.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\0n0wze2r.g2o","hash":"mx+2/l60CP8o8HN/ojT+PQ=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"client-alert-notifications-by-email\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/get-started/alert-email-notifications.md\" sourcestartlinenumber=\"25\">Client-Warnungsbenachrichtigungen per E-Mail</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/02_SupportProcesses/02_03_Project/Project2.md","output":{".html":{"relative_path":"ProcessDoku/02_SupportProcesses/02_03_Project/Project2.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\q2kullhh.mzh","hash":"qBRMsi19+5SOmcs/TLDv9g=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"ProcessDoku/01_CoreProcesses/01_09_Invoicing/Invoicing.md","output":{".html":{"relative_path":"ProcessDoku/01_CoreProcesses/01_09_Invoicing/Invoicing.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\sodpw1mm.aiy","hash":"YZKCM2aBdqxJwLodnIsVfw=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"invoicing\" sourcefile=\"ProcessDoku/01_CoreProcesses/01_09_Invoicing/Invoicing.md\" sourcestartlinenumber=\"1\">Invoicing</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/01_CoreProcesses/01_08_Receiving/Receiving2.md","output":{".html":{"relative_path":"ProcessDoku/01_CoreProcesses/01_08_Receiving/Receiving2.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\mcrlov0k.xix","hash":"wybnbxCAJGo8z0m3l4l5mQ=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"receiving-2\" sourcefile=\"ProcessDoku/01_CoreProcesses/01_08_Receiving/Receiving2.md\" sourcestartlinenumber=\"1\">Receiving 2</h1>"},{"log_codes":["InvalidFileLink"],"type":"Conceptual","source_relative_path":"ProcessDoku/01_CoreProcesses/01_04_Production/Production.md","output":{".html":{"relative_path":"ProcessDoku/01_CoreProcesses/01_04_Production/Production.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\buf2atsv.nwz","hash":"G3kng0Z6AhGCbp6b84h5/Q=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"production-process-overview\" sourcefile=\"ProcessDoku/01_CoreProcesses/01_04_Production/Production.md\" sourcestartlinenumber=\"5\">Production process overview</h1>"},{"log_codes":["InvalidFileLink"],"type":"Conceptual","source_relative_path":"ProcessDoku/01_CoreProcesses/01_04_Production/ProdPlanning_Overview.md","output":{".html":{"relative_path":"ProcessDoku/01_CoreProcesses/01_04_Production/ProdPlanning_Overview.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\mcyjxryr.cfh","hash":"VARqqzt9hPfBA5fiAWxebw=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"production-planning\" sourcefile=\"ProcessDoku/01_CoreProcesses/01_04_Production/ProdPlanning_Overview.md\" sourcestartlinenumber=\"1\">PRODUCTION PLANNING</h1>"},{"log_codes":["InvalidFileLink"],"type":"Conceptual","source_relative_path":"ProcessDoku/01_CoreProcesses/01_01_CRM/CRM2.md","output":{".html":{"relative_path":"ProcessDoku/01_CoreProcesses/01_01_CRM/CRM2.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\lyfzsxbu.hyx","hash":"xODoRGd1OASCQaiMAcVxIA=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"crm2\" sourcefile=\"ProcessDoku/01_CoreProcesses/01_01_CRM/CRM2.md\" sourcestartlinenumber=\"1\">CRM2</h1>"},{"log_codes":["InvalidFileLink"],"type":"Conceptual","source_relative_path":"ProcessDoku/01_CoreProcesses/01_01_CRM/CRM1.md","output":{".html":{"relative_path":"ProcessDoku/01_CoreProcesses/01_01_CRM/CRM1.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\4hbm3i3r.dwa","hash":"P2kHugvmgomV+6RGSEWfBg=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"crm\" sourcefile=\"ProcessDoku/01_CoreProcesses/01_01_CRM/CRM1.md\" sourcestartlinenumber=\"1\">CRM</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/set-up-number-sequences-individual-basis.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/set-up-number-sequences-individual-basis.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\ftkextcc.ykj","hash":"8GLvgGvOUw64ispRkQGoJA=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"set-up-number-sequences-on-an-individual-basis\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/set-up-number-sequences-individual-basis.md\" sourcestartlinenumber=\"25\">Nummernkreise einzeln einrichten</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/set-up-electronic-signatures.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/set-up-electronic-signatures.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\3eqzjest.m5c","hash":"LcK726b+e6iYKxdQQZTzIA=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"set-up-electronic-signatures\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/set-up-electronic-signatures.md\" sourcestartlinenumber=\"25\">Einrichten elektronischer Signaturen</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/workflow-actions.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/workflow-actions.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\upiyihpj.u5g","hash":"QGD0AiSILamTvnocaa4lXw=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"actions-in-workflow-approval-processes\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/organization-administration/workflow-actions.md\" sourcestartlinenumber=\"26\">Aktivitäten in Workflow-Genehmigungsprozessen</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/record-templates.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/record-templates.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\3lysrklg.q54","hash":"yiz2ZkkEWA7abUoIuEycUw=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"record-templates-overview\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/organization-administration/record-templates.md\" sourcestartlinenumber=\"26\">Übersicht über die Aufnahmevorlagen</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/number-sequence-overview.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/number-sequence-overview.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\kldqiiaa.nro","hash":"pQRJsS3Mbh2PSX7W/R71kQ=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"number-sequences-overview\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/organization-administration/number-sequence-overview.md\" sourcestartlinenumber=\"27\">Nummernkreisübersicht</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/electronic-signature-overview.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/electronic-signature-overview.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\rewwdu5e.lg2","hash":"He/I67KV8tk9N8uyD/Sqmw=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"electronic-signatures-overview\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/organization-administration/electronic-signature-overview.md\" sourcestartlinenumber=\"27\">Elektronische Signatur – Übersicht</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/configure-manual-task-workflow.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/configure-manual-task-workflow.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\nzsg02je.ov3","hash":"+dNHt08bXweZgZIqHDDHIg=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"configure-manual-tasks-in-a-workflow\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/organization-administration/configure-manual-task-workflow.md\" sourcestartlinenumber=\"26\">Manuelle Aufgaben in einem Workflow konfigurieren</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/hr/tasks/manage-leave-absence.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/hr/tasks/manage-leave-absence.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\s4kvgsfq.ill","hash":"gTGOJjVbxG8Sm/np7VHcrg=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"manage-leave-of-absence\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/hr/tasks/manage-leave-absence.md\" sourcestartlinenumber=\"25\">Beurlaubung verwalten</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/hr/tasks/approve-application-inbox-records.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/hr/tasks/approve-application-inbox-records.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\hspn4off.a4d","hash":"ZeDIQRKfhJey6TfzIuCMmA=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"approve-application-inbox-records\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/hr/tasks/approve-application-inbox-records.md\" sourcestartlinenumber=\"25\">Bewerbungseingangs-Datensätze genehmigen</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/01_CoreProcesses/01_05_Purchasing/Purchasing2.md","output":{".html":{"relative_path":"ProcessDoku/01_CoreProcesses/01_05_Purchasing/Purchasing2.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\yvbpx2gt.lhz","hash":"pzOYgPpjG16NOAHivxaasg=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"purchasing-2\" sourcefile=\"ProcessDoku/01_CoreProcesses/01_05_Purchasing/Purchasing2.md\" sourcestartlinenumber=\"1\">Purchasing 2</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/01_CoreProcesses/01_05_Purchasing/Purchasing1.md","output":{".html":{"relative_path":"ProcessDoku/01_CoreProcesses/01_05_Purchasing/Purchasing1.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\fnfyjbkm.p45","hash":"Xi5n8kpLri6CtDFoOchRrQ=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"purchasing-1\" sourcefile=\"ProcessDoku/01_CoreProcesses/01_05_Purchasing/Purchasing1.md\" sourcestartlinenumber=\"1\">Purchasing 1</h1>"},{"log_codes":["include-not-found"],"type":"Conceptual","source_relative_path":"ProcessDoku/01_CoreProcesses/01_02_Quotations/Quotations2.md","output":{".html":{"relative_path":"ProcessDoku/01_CoreProcesses/01_02_Quotations/Quotations2.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\2qmnzqvo.5qy","hash":"mqov71jsNej6HUlWJiB6JA=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"price-simulation\" sourcefile=\"ProcessDoku/01_CoreProcesses/01_02_Quotations/Quotations2.md\" sourcestartlinenumber=\"1\">Price simulation</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/view-workflow-history.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/view-workflow-history.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\f0hj5e4w.fr3","hash":"Wuu0PiGLZrkVOoj01GjbHg=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"view-workflow-history\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/view-workflow-history.md\" sourcestartlinenumber=\"25\">Anzeigen der Workflowhistorie</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/users-receive-workflow-related-email-messages.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/users-receive-workflow-related-email-messages.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\aps14tsz.td2","hash":"hYUKruSLqvv68nEkdFBc8w=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"enable-users-to-receive-workflow-related-email-messages\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/users-receive-workflow-related-email-messages.md\" sourcestartlinenumber=\"25\">Ermöglichen Sie es Benutzern, workflowbezogene E-Mail-Nachrichten zu erhalten.</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/create-operating-unit.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/create-operating-unit.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\3apekdg5.j0p","hash":"KA1RsnceqlAcFhzFWeUYwA=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"create-an-operating-unit\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/create-operating-unit.md\" sourcestartlinenumber=\"25\">Organisationseinheit erstellen</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/includes/preview-banner.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/includes/preview-banner.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\tp2qa1lw.ak5","hash":"ZlVEZJ4KEFyY3i9HSJ6WFw=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/hr/tasks/identify-deploy-candidate-selection-tools.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/hr/tasks/identify-deploy-candidate-selection-tools.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\rovewftc.xda","hash":"YzY+CY+0b1LgenBul4jLbQ=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"identify-and-deploy-candidate-selection-tools\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/hr/tasks/identify-deploy-candidate-selection-tools.md\" sourcestartlinenumber=\"25\">Hilfsmittel zur Kandidatenauswahl ermitteln und bereitstellen</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/hr/localizations/noam-usa-enter-beginning-balances.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/hr/localizations/noam-usa-enter-beginning-balances.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\hq0ilq3t.gwr","hash":"zF3twOaOIsuaRJ4WL7G7EA=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"enter-payroll-beginning-balances\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/hr/localizations/noam-usa-enter-beginning-balances.md\" sourcestartlinenumber=\"26\">Eingeben von Lohnanfangssalden</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/user-interface-elements.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/user-interface-elements.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\dhay3r35.zm4","hash":"Wiytle0ADYb4YvxQvTmTMg=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"user-interface-elements\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/get-started/user-interface-elements.md\" sourcestartlinenumber=\"24\">Benutzeroberflächenelemente</h1>"},{"log_codes":["include-not-found"],"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/change-date-session.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/change-date-session.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\ehmyv4bl.zmg","hash":"nQZP7yPfCLqHg2cONtFo/g=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"change-the-date-for-a-session\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/get-started/change-date-session.md\" sourcestartlinenumber=\"25\">Ändern des Datums für eine Sitzung</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/accessibility-features.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/accessibility-features.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\ozvihdzk.tkh","hash":"8Q/58i5YNJ7oEPLlXpBK2g=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"accessibility-features\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/get-started/accessibility-features.md\" sourcestartlinenumber=\"24\">Eingabehilfefunktionen</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/03_GlobalDataAndDataExchange/03_03_GDDS/GDDS2.md","output":{".html":{"relative_path":"ProcessDoku/03_GlobalDataAndDataExchange/03_03_GDDS/GDDS2.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\n5r30vxz.0jf","hash":"Mt9SmE/f9Wz0Pvi/xf+eIA=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"ProcessDoku/03_GlobalDataAndDataExchange/03_03_GDDS/GDDS1.md","output":{".html":{"relative_path":"ProcessDoku/03_GlobalDataAndDataExchange/03_03_GDDS/GDDS1.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\eesmgitc.yuh","hash":"rwvolN1AvcAwsqLxos9yBw=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"ProcessDoku/02_SupportProcesses/02_03_Project/Project_Overview.md","output":{".html":{"relative_path":"ProcessDoku/02_SupportProcesses/02_03_Project/Project_Overview.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\lfckjudc.400","hash":"517KJQc7/kD8m9srq4u0sg=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"ProcessDoku/03_GlobalDataAndDataExchange/GdAndDe_Overview.md","output":{".html":{"relative_path":"ProcessDoku/03_GlobalDataAndDataExchange/GdAndDe_Overview.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\t12j4bsz.dtw","hash":"mHe2zumlreuU0H1UAT2jCg=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"global-data-and-data-exchange-overview\" sourcefile=\"ProcessDoku/03_GlobalDataAndDataExchange/GdAndDe_Overview.md\" sourcestartlinenumber=\"1\">Global Data and Data Exchange Overview</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/02_SupportProcesses/02_04_ECN/ECN_Overview.md","output":{".html":{"relative_path":"ProcessDoku/02_SupportProcesses/02_04_ECN/ECN_Overview.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\tbopbwib.zqv","hash":"28QGF2t7iggtRnwcV4lQcw=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"ProcessDoku/03_GlobalDataAndDataExchange/03_01_RemoteCall/RemoteCall_Overview.md","output":{".html":{"relative_path":"ProcessDoku/03_GlobalDataAndDataExchange/03_01_RemoteCall/RemoteCall_Overview.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\fnu0hocw.kto","hash":"Lkr179AyOMAtQZaulN91Eg=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"ProcessDoku/02_SupportProcesses/02_02_ServiceProcesses/02_02_01_Maintenance/Maintenance1.md","output":{".html":{"relative_path":"ProcessDoku/02_SupportProcesses/02_02_ServiceProcesses/02_02_01_Maintenance/Maintenance1.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\oo1uiila.nle","hash":"y8SqOATj0vTEjw8de1RZOA=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"ProcessDoku/02_SupportProcesses/02_02_ServiceProcesses/ServiceProcesses_Overview.md","output":{".html":{"relative_path":"ProcessDoku/02_SupportProcesses/02_02_ServiceProcesses/ServiceProcesses_Overview.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\1snawpqy.xpc","hash":"nAjL8wOtNvuMj7GF8jlLvQ=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"ProcessDoku/02_SupportProcesses/SupportProcesses_Overview.md","output":{".html":{"relative_path":"ProcessDoku/02_SupportProcesses/SupportProcesses_Overview.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\oy5odu0j.ukb","hash":"UH1t/Rm49OHG0Sgx1yR74Q=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"support-processes-overview\" sourcefile=\"ProcessDoku/02_SupportProcesses/SupportProcesses_Overview.md\" sourcestartlinenumber=\"1\">Support Processes Overview</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/01_CoreProcesses/01_10_ModelcodeGuideline/ModelcodeGuideline2.md","output":{".html":{"relative_path":"ProcessDoku/01_CoreProcesses/01_10_ModelcodeGuideline/ModelcodeGuideline2.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\g3wtobkr.bij","hash":"ewxZz1e4Z9L1o2i4n1nNYg=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"modelcodeguideline2\" sourcefile=\"ProcessDoku/01_CoreProcesses/01_10_ModelcodeGuideline/ModelcodeGuideline2.md\" sourcestartlinenumber=\"1\">ModelcodeGuideline2</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/01_CoreProcesses/01_06_Warehouse/Warehouse1.md","output":{".html":{"relative_path":"ProcessDoku/01_CoreProcesses/01_06_Warehouse/Warehouse1.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\jxnwtvwu.vqc","hash":"kvq4DUU4rlekJ7wHaUU4IA=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"warehouse-1\" sourcefile=\"ProcessDoku/01_CoreProcesses/01_06_Warehouse/Warehouse1.md\" sourcestartlinenumber=\"1\">Warehouse 1</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/02_SupportProcesses/02_01_Finance/Finance2.md","output":{".html":{"relative_path":"ProcessDoku/02_SupportProcesses/02_01_Finance/Finance2.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\twduqtsx.s4u","hash":"ZnjKBK8mg0xswEvoMJrQXQ=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"ProcessDoku/02_SupportProcesses/02_01_Finance/Finance1.md","output":{".html":{"relative_path":"ProcessDoku/02_SupportProcesses/02_01_Finance/Finance1.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\aw0gnu5k.zhj","hash":"VZaCO7T476VjSON5DElF9Q=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"ProcessDoku/01_CoreProcesses/01_08_Receiving/Receiving1.md","output":{".html":{"relative_path":"ProcessDoku/01_CoreProcesses/01_08_Receiving/Receiving1.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\dojhkglf.fkn","hash":"Wh5n4mkbiDme61+A4L9mIg=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"receiving-1\" sourcefile=\"ProcessDoku/01_CoreProcesses/01_08_Receiving/Receiving1.md\" sourcestartlinenumber=\"1\">Receiving 1</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/01_CoreProcesses/01_08_Receiving/Receiving.md","output":{".html":{"relative_path":"ProcessDoku/01_CoreProcesses/01_08_Receiving/Receiving.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\f2ovhjaa.g1h","hash":"LzEBuUt2gyDQq0iKGXdlKg=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"receiving\" sourcefile=\"ProcessDoku/01_CoreProcesses/01_08_Receiving/Receiving.md\" sourcestartlinenumber=\"1\">Receiving</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/01_CoreProcesses/01_06_Warehouse/Warehouse.md","output":{".html":{"relative_path":"ProcessDoku/01_CoreProcesses/01_06_Warehouse/Warehouse.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\ewcnx5tn.dtf","hash":"FkUqgC0soWAxoTG+ZDaNQQ=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"warehouse\" sourcefile=\"ProcessDoku/01_CoreProcesses/01_06_Warehouse/Warehouse.md\" sourcestartlinenumber=\"1\">Warehouse</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/01_CoreProcesses/01_03_Sales/Sales_Agreements.md","output":{".html":{"relative_path":"ProcessDoku/01_CoreProcesses/01_03_Sales/Sales_Agreements.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\1wvlivac.mld","hash":"HtrTKGuvxigZYKgMAZ18qw=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"sales-agreements-overview\" sourcefile=\"ProcessDoku/01_CoreProcesses/01_03_Sales/Sales_Agreements.md\" sourcestartlinenumber=\"5\">Sales agreements overview</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/set-users-preferred-time-zone.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/set-users-preferred-time-zone.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\rfvrvu4x.eqc","hash":"cZZQd5iptMUCnWNPAxjQ0A=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"set-a-users-preferred-time-zone\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/set-users-preferred-time-zone.md\" sourcestartlinenumber=\"25\">Die bevorzugte Zeitzone eines Benutzers festlegen</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/set-up-number-sequences-wizard.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/set-up-number-sequences-wizard.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\vzbfbs0f.hd2","hash":"pOyjr+Lf8HkmjsTR43n1Hg=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"set-up-number-sequences-using-a-wizard\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/set-up-number-sequences-wizard.md\" sourcestartlinenumber=\"25\">Einrichten von Nummernkreisen mit einem Assistenten</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/change-date-session.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/change-date-session.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\xmbrr05n.23e","hash":"ArY4+kbO+dzD+BtKb64vcg=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"change-the-date-for-a-session\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/change-date-session.md\" sourcestartlinenumber=\"25\">Ändern des Datums für eine Sitzung</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/address-books.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/address-books.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\v54my4gh.ie2","hash":"ABPolil7vvYpHPdvzDcKEw=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"configure-address-books\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/address-books.md\" sourcestartlinenumber=\"25\">Adressbücher konfigurieren</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/create-workflow.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/create-workflow.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\mournjtu.ns4","hash":"t1QsYHo1VqVj625fE9Uxhw=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"create-workflows-overview\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/organization-administration/create-workflow.md\" sourcestartlinenumber=\"27\">Erstellen von Workflows – Übersicht</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/configure-workflow-properties.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/configure-workflow-properties.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\jgrbxogm.qdy","hash":"MiOUlYTtB64ScUp4pwQczg=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"configure-workflow-properties\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/organization-administration/configure-workflow-properties.md\" sourcestartlinenumber=\"26\">Konfigurieren von Workfloweigenschaften</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/hr/tasks/enter-applicant-application-data-manually.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/hr/tasks/enter-applicant-application-data-manually.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\5mpdtnc1.nou","hash":"PtCQUO9yBBf4Q6RuFh03TA=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"enter-applicant-and-application-data-manually\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/hr/tasks/enter-applicant-application-data-manually.md\" sourcestartlinenumber=\"25\">Bewerber- und Anwendungsdaten manuell eingeben</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/hr/tasks/develop-open-job-requisition.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/hr/tasks/develop-open-job-requisition.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\vu2scm1w.1kx","hash":"nndnOH/VvL+cx/8Xao7k9w=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"develop-and-open-job-requisition\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/hr/tasks/develop-open-job-requisition.md\" sourcestartlinenumber=\"25\">Stellenanforderung ausarbeiten und freigeben</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/tasks/change-banner-or-logo.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/tasks/change-banner-or-logo.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\f1vjyuvn.4uy","hash":"PpOz83xJue3ADp1bU5J/yA=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"change-the-banner-or-logo\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/get-started/tasks/change-banner-or-logo.md\" sourcestartlinenumber=\"25\">Das Banner oder das Logo ändern</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/action-search.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/action-search.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\jqqutm3z.4wf","hash":"adU6CBLXUtFMxTESiAcNRg=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"action-search\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/get-started/action-search.md\" sourcestartlinenumber=\"26\">Aktivitätssuche</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/02_SupportProcesses/02_03_Project/Project1.md","output":{".html":{"relative_path":"ProcessDoku/02_SupportProcesses/02_03_Project/Project1.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\yl4ir4km.njt","hash":"Lj3xsSgOpB/2uuitinc0Rw=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"ProcessDoku/02_SupportProcesses/02_04_ECN/ECN2.md","output":{".html":{"relative_path":"ProcessDoku/02_SupportProcesses/02_04_ECN/ECN2.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\yu3k1yuw.4u2","hash":"0Mt6hGn2eejFXBtxXT3tiQ=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"ProcessDoku/02_SupportProcesses/02_04_ECN/ECN1.md","output":{".html":{"relative_path":"ProcessDoku/02_SupportProcesses/02_04_ECN/ECN1.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\ojkumcwe.ecz","hash":"V727Ain0WJIKrNPe6cHtTQ=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"ProcessDoku/02_SupportProcesses/02_02_ServiceProcesses/02_02_01_Maintenance/Maintenance_Overview.md","output":{".html":{"relative_path":"ProcessDoku/02_SupportProcesses/02_02_ServiceProcesses/02_02_01_Maintenance/Maintenance_Overview.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\i4nh3ijw.px4","hash":"iDg0rCGo0+ssqZogxnB/UA=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"ProcessDoku/02_SupportProcesses/02_02_ServiceProcesses/02_02_01_Maintenance/Maintenance2.md","output":{".html":{"relative_path":"ProcessDoku/02_SupportProcesses/02_02_ServiceProcesses/02_02_01_Maintenance/Maintenance2.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\zof2k3ba.utv","hash":"BMV3JM6RYWkj1h98XxSOuQ=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"ProcessDoku/01_CoreProcesses/01_09_Invoicing/Invoicing2.md","output":{".html":{"relative_path":"ProcessDoku/01_CoreProcesses/01_09_Invoicing/Invoicing2.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\mhkqrrkh.gt2","hash":"k3Sa25abyHzJDfPtEnIzuQ=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"invoicing-2\" sourcefile=\"ProcessDoku/01_CoreProcesses/01_09_Invoicing/Invoicing2.md\" sourcestartlinenumber=\"1\">Invoicing 2</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/01_CoreProcesses/01_09_Invoicing/Invoicing1.md","output":{".html":{"relative_path":"ProcessDoku/01_CoreProcesses/01_09_Invoicing/Invoicing1.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\pfbjmqbt.pfg","hash":"Tr2fb/y+2vXWSXXZTGMfzA=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"invoicing-1\" sourcefile=\"ProcessDoku/01_CoreProcesses/01_09_Invoicing/Invoicing1.md\" sourcestartlinenumber=\"1\">Invoicing 1</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/01_CoreProcesses/01_07_Shipping/Shipping.md","output":{".html":{"relative_path":"ProcessDoku/01_CoreProcesses/01_07_Shipping/Shipping.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\vm5twllp.rfy","hash":"dpNS8ca9EiktTF2xLCuseQ=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"shipping\" sourcefile=\"ProcessDoku/01_CoreProcesses/01_07_Shipping/Shipping.md\" sourcestartlinenumber=\"1\">Shipping</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/01_CoreProcesses/01_06_Warehouse/Warehouse2.md","output":{".html":{"relative_path":"ProcessDoku/01_CoreProcesses/01_06_Warehouse/Warehouse2.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\e4en0vtm.lsq","hash":"mT4bEEpuGPgjVU7I+Z6jMA=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"warehouse-2\" sourcefile=\"ProcessDoku/01_CoreProcesses/01_06_Warehouse/Warehouse2.md\" sourcestartlinenumber=\"1\">Warehouse 2</h1>"},{"log_codes":["InvalidFileLink"],"type":"Conceptual","source_relative_path":"ProcessDoku/01_CoreProcesses/01_04_Production/ProdPlanning2.md","output":{".html":{"relative_path":"ProcessDoku/01_CoreProcesses/01_04_Production/ProdPlanning2.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\ae3e2fdy.g5y","hash":"3Gt9jomdCW6Msp2VEEQiBw=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"production-planning-2\" sourcefile=\"ProcessDoku/01_CoreProcesses/01_04_Production/ProdPlanning2.md\" sourcestartlinenumber=\"1\">Production Planning 2</h1>"},{"log_codes":["InvalidFileLink"],"type":"Conceptual","source_relative_path":"ProcessDoku/01_CoreProcesses/01_04_Production/ProdPlanning1.md","output":{".html":{"relative_path":"ProcessDoku/01_CoreProcesses/01_04_Production/ProdPlanning1.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\gsygzpsm.cx2","hash":"9Sgtf8x24MIr6Le7MpiN+A=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"production-planning-1\" sourcefile=\"ProcessDoku/01_CoreProcesses/01_04_Production/ProdPlanning1.md\" sourcestartlinenumber=\"1\">Production Planning 1</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/01_CoreProcesses/01_02_Quotations/Quotations1.md","output":{".html":{"relative_path":"ProcessDoku/01_CoreProcesses/01_02_Quotations/Quotations1.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\suyszhcu.to2","hash":"LxO7ICner1cFWfUIi0TF0w=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"mass-create-sales-quotations\" sourcefile=\"ProcessDoku/01_CoreProcesses/01_02_Quotations/Quotations1.md\" sourcestartlinenumber=\"1\">Mass create sales quotations</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/delegate-work-items-workflow.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/delegate-work-items-workflow.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\ff22mmab.lqd","hash":"Hl/kRv+/TwIxjbgcvXjbzw=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"delegate-work-items-in-a-workflow\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/delegate-work-items-workflow.md\" sourcestartlinenumber=\"25\">Delegieren von Arbeitsaufgaben in einem Workflow</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/create-organization-hierarchy.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/create-organization-hierarchy.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\me4tvep3.rkc","hash":"3XGjdID86y0Kn571bw7Z2Q=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"create-an-organization-hierarchy\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/organization-administration/tasks/create-organization-hierarchy.md\" sourcestartlinenumber=\"25\">Erstellen Sie eine Organisationshierarchie</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/workflow-FAQ.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/workflow-FAQ.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\bdflund2.es0","hash":"AUhQHnrmMs6x9IEYK3saeA=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"workflow-faq\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/organization-administration/workflow-FAQ.md\" sourcestartlinenumber=\"24\">Workflow-FAQs</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/workflow-elements.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/workflow-elements.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\r3h2uzec.f2k","hash":"CJMUqMTgWcyXg4jNWNUL0A=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"workflow-elements\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/organization-administration/workflow-elements.md\" sourcestartlinenumber=\"26\">Workflowelemente</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/shortcut-keys.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/shortcut-keys.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\va5zjdbt.b3n","hash":"2USyiHeRQ7wroajxH/kfOw=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"keyboard-shortcuts\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/get-started/shortcut-keys.md\" sourcestartlinenumber=\"26\">Tastenkombinationen</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/navigation-search.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/navigation-search.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\thw35vf4.miz","hash":"epIfmbsAZjXa8vsu6R2C6Q=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"navigation-search\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/get-started/navigation-search.md\" sourcestartlinenumber=\"26\">Navigationssuche</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/alerts-overview.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/alerts-overview.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\15znmtd1.3f5","hash":"Gq2TyPk/y+fNyYFgjtMZ0A=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"alerts-overview\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/get-started/alerts-overview.md\" sourcestartlinenumber=\"25\">Überblick über Warnungen</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/advanced-filtering-query-options.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/advanced-filtering-query-options.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\1kf0ybzt.cg1","hash":"meEAZERUpqjEsouIelIm4A=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"advanced-filtering-and-query-syntax\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/get-started/advanced-filtering-query-options.md\" sourcestartlinenumber=\"27\">Erweiterte Filter- und Abfragesyntax</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/Notifications.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/Notifications.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\hj0f4zje.p4o","hash":"lW7RRzkpYJi726KvRIs3IQ=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"what-exactly-are-notifications\" sourcefile=\"ProcessDoku/00_Basics/Notifications.md\" sourcestartlinenumber=\"1\">WHAT EXACTLY ARE NOTIFICATIONS</h1>"},{"log_codes":["InvalidFileLink"],"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/Login.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/Login.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\p3wqph3o.t3h","hash":"lGvqfQXj462l7eGhUhltDQ=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"login\" sourcefile=\"ProcessDoku/00_Basics/Login.md\" sourcestartlinenumber=\"1\">Login</h1>"},{"log_codes":["InvalidFileLink"],"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/Basics.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/Basics.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\h35byjhp.m3n","hash":"iM3zc07MBVLYzXlMEa0q0A=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"basics\" sourcefile=\"ProcessDoku/00_Basics/Basics.md\" sourcestartlinenumber=\"1\">Basics</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/03_GlobalDataAndDataExchange/03_03_GDDS/GDDS_Overview.md","output":{".html":{"relative_path":"ProcessDoku/03_GlobalDataAndDataExchange/03_03_GDDS/GDDS_Overview.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\dtz3s54n.hdq","hash":"mZwZdp4vTPSjqTC2irCwvA=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"ProcessDoku/02_SupportProcesses/02_02_ServiceProcesses/02_02_02_InstalledBase/InstalledBase2.md","output":{".html":{"relative_path":"ProcessDoku/02_SupportProcesses/02_02_ServiceProcesses/02_02_02_InstalledBase/InstalledBase2.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\zkdrkknp.h5j","hash":"bXhFW/tBTIaAz8WZyk3B0A=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"ProcessDoku/02_SupportProcesses/02_02_ServiceProcesses/02_02_02_InstalledBase/InstalledBase1.md","output":{".html":{"relative_path":"ProcessDoku/02_SupportProcesses/02_02_ServiceProcesses/02_02_02_InstalledBase/InstalledBase1.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\u2h4qa3v.wrv","hash":"Xfj7k6uhKp+WKTWDsCnTFQ=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"ProcessDoku/01_CoreProcesses/01_07_Shipping/Shipping2.md","output":{".html":{"relative_path":"ProcessDoku/01_CoreProcesses/01_07_Shipping/Shipping2.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\ed124lot.z14","hash":"i7cAH1bP+QqhvMf7wB4d6Q=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"shipping-2\" sourcefile=\"ProcessDoku/01_CoreProcesses/01_07_Shipping/Shipping2.md\" sourcestartlinenumber=\"1\">Shipping 2</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/01_CoreProcesses/01_07_Shipping/Shipping1.md","output":{".html":{"relative_path":"ProcessDoku/01_CoreProcesses/01_07_Shipping/Shipping1.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\2kwokwus.0hk","hash":"yEy3wm6hk5tTszrFpjd2PQ=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"shipping-1\" sourcefile=\"ProcessDoku/01_CoreProcesses/01_07_Shipping/Shipping1.md\" sourcestartlinenumber=\"1\">Shipping 1</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/01_CoreProcesses/01_05_Purchasing/Purchasing.md","output":{".html":{"relative_path":"ProcessDoku/01_CoreProcesses/01_05_Purchasing/Purchasing.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\al3p0wcm.rnj","hash":"fuIkV8cW5kbwgdRcSFsypw=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"add-your-introductions-here\" sourcefile=\"ProcessDoku/01_CoreProcesses/01_05_Purchasing/Purchasing.md\" sourcestartlinenumber=\"1\">Add your introductions here!</h1>"},{"log_codes":["InvalidFileLink"],"type":"Conceptual","source_relative_path":"ProcessDoku/01_CoreProcesses/01_04_Production/PROD_Ressoucen.md","output":{".html":{"relative_path":"ProcessDoku/01_CoreProcesses/01_04_Production/PROD_Ressoucen.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\j3smmmvp.bug","hash":"IucZBWKZ0hc4XAq7gj99LQ=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"ressourcen-in-d365\" sourcefile=\"ProcessDoku/01_CoreProcesses/01_04_Production/PROD_Ressoucen.md\" sourcestartlinenumber=\"2\">Ressourcen in D365</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/02_SupportProcesses/02_02_ServiceProcesses/02_02_02_InstalledBase/InstalledBase_Overview.md","output":{".html":{"relative_path":"ProcessDoku/02_SupportProcesses/02_02_ServiceProcesses/02_02_02_InstalledBase/InstalledBase_Overview.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\cbzu23xs.nww","hash":"91ukSp2UpBB7nlYYDXVg7w=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/organizations-organizational-hierarchies.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/organizations-organizational-hierarchies.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\i14u551v.hgn","hash":"/EIDwhv0VHZ8lZYJFElG2A=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"organizations-and-organizational-hierarchies-overview\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/organization-administration/organizations-organizational-hierarchies.md\" sourcestartlinenumber=\"27\">Übersicht über Unternehmen und Organisationshierarchien</h1>"},{"log_codes":["InvalidFileLink"],"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/organization-administration-home-page.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/organization-administration-home-page.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\czo25vq1.ufc","hash":"AcAt8ccGgvctfNLMVUrE0A=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"organization-administration-home-page\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/organization-administration/organization-administration-home-page.md\" sourcestartlinenumber=\"26\">Organisationsverwaltung – Startseite</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/configure-approval-process-workflow.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/configure-approval-process-workflow.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\aazisjx4.pi4","hash":"f3z7dHPSiWYPaElnDZQ1jQ=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"configure-approval-processes-in-a-workflow\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/organization-administration/configure-approval-process-workflow.md\" sourcestartlinenumber=\"26\">Genehmigungsprozesse in einem Workflow konfigurieren</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/includes/banner.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/includes/banner.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\lq1sah5n.fkw","hash":"jaT5jqWKV58AgGtlUsGASw=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/hr/tasks/hire-existing-employee-through-recruiting.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/hr/tasks/hire-existing-employee-through-recruiting.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\nhtpyaab.ghg","hash":"sxZFYL96d5OY/qo3LxiMHw=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"hire-existing-employees-through-recruitment\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/hr/tasks/hire-existing-employee-through-recruiting.md\" sourcestartlinenumber=\"24\">Vorhandene Mitarbeiter mittels Personalbeschaffung einstellen</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/hr/manage-recruiting-process.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/hr/manage-recruiting-process.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\hd2zvq4o.d1e","hash":"IgVgJJVLm0CYjUG4SX0ZKA=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"manage-recruiting-processes\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/hr/manage-recruiting-process.md\" sourcestartlinenumber=\"27\">Personalbeschaffungsprozesse verwalten</h1>"},{"log_codes":["include-not-found"],"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/set-users-preferred-time-zone.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/set-users-preferred-time-zone.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\eho1kwbm.343","hash":"kaPRiPWix5DMw4p4Wi/M2w=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"set-a-users-preferred-time-zone\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/get-started/set-users-preferred-time-zone.md\" sourcestartlinenumber=\"25\">Die bevorzugte Zeitzone eines Benutzers festlegen</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/display-pages-side-by-side.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/display-pages-side-by-side.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\3mqtvod2.3pr","hash":"0ZlIKz18yYO16G4WE3OOOQ=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"show-pages-side-by-side-using-the-open-in-new-window-feature\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/get-started/display-pages-side-by-side.md\" sourcestartlinenumber=\"26\">Seiten mithilfe der Funktion „In neuem Fenster öffnen“ nebeneinander anzeigen</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/alerts-managing.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/alerts-managing.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\agno41yi.b2u","hash":"NihoPRW2CLdlhvx3p7MSjA=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"batch-processing-of-alerts\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/get-started/alerts-managing.md\" sourcestartlinenumber=\"24\">Stapelverarbeitung von Warnungen</h1>"},{"log_codes":["InvalidFileLink"],"type":"Conceptual","source_relative_path":"ProcessDoku/intro.md","output":{".html":{"relative_path":"ProcessDoku/intro.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\413mgulj.4gp","hash":"7wG2V+zdxHS59yQrIHwktA=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"welcome-page-wika-process-doku\" sourcefile=\"ProcessDoku/intro.md\" sourcestartlinenumber=\"1\">Welcome Page WIKA Process Doku</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/03_GlobalDataAndDataExchange/03_01_RemoteCall/RemoteCall2.md","output":{".html":{"relative_path":"ProcessDoku/03_GlobalDataAndDataExchange/03_01_RemoteCall/RemoteCall2.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\t0sl2hrf.ixg","hash":"XhJSQuTWhT6iaMgEGPJmag=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"ProcessDoku/03_GlobalDataAndDataExchange/03_01_RemoteCall/RemoteCall1.md","output":{".html":{"relative_path":"ProcessDoku/03_GlobalDataAndDataExchange/03_01_RemoteCall/RemoteCall1.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\n5nojwui.cwj","hash":"/xFtKHnxa/y+eNezJ3g1bQ=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"ProcessDoku/02_SupportProcesses/02_02_ServiceProcesses/ServiceProcesses1.md","output":{".html":{"relative_path":"ProcessDoku/02_SupportProcesses/02_02_ServiceProcesses/ServiceProcesses1.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\bf3qk1hv.mmb","hash":"NHqC08z2M6xjdJM1BU8wyw=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"ProcessDoku/02_SupportProcesses/02_01_Finance/Finance_Overview.md","output":{".html":{"relative_path":"ProcessDoku/02_SupportProcesses/02_01_Finance/Finance_Overview.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\b120qptp.e2x","hash":"ytRt52WdP3A4LhoDJ7+x/w=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"ProcessDoku/01_CoreProcesses/01_10_ModelcodeGuideline/ModelcodeGuideline1.md","output":{".html":{"relative_path":"ProcessDoku/01_CoreProcesses/01_10_ModelcodeGuideline/ModelcodeGuideline1.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\5cddxipi.pnv","hash":"41V+iFBAboRJovcVs18XuQ=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"modelcodeguideline1\" sourcefile=\"ProcessDoku/01_CoreProcesses/01_10_ModelcodeGuideline/ModelcodeGuideline1.md\" sourcestartlinenumber=\"1\">ModelcodeGuideline1</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/01_CoreProcesses/01_10_ModelcodeGuideline/ModelcodeGuideline.md","output":{".html":{"relative_path":"ProcessDoku/01_CoreProcesses/01_10_ModelcodeGuideline/ModelcodeGuideline.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\44tmwakm.5dt","hash":"UHdhAMMIPzcGkp40/spPOg=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"modelcodeguideline\" sourcefile=\"ProcessDoku/01_CoreProcesses/01_10_ModelcodeGuideline/ModelcodeGuideline.md\" sourcestartlinenumber=\"1\">ModelcodeGuideline</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/plan-configuration-global-address-book-additional-address-books.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/plan-configuration-global-address-book-additional-address-books.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\0h0uspsc.nhw","hash":"CmpGNWJ3nb/8iXZT/UVvCg=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"plan-for-the-global-address-book-and-other-address-books\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/organization-administration/plan-configuration-global-address-book-additional-address-books.md\" sourcestartlinenumber=\"27\">Planen für das globale Adressbuch und andere Adressbücher</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/overview-workflow-system.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/overview-workflow-system.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\lkpdhz3p.wtt","hash":"YYVihH07o/TO/n4qtOZ/Zw=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"workflow-system-overview\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/organization-administration/overview-workflow-system.md\" sourcestartlinenumber=\"26\">Workflowsystem – Übersicht</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/configure-line-item-workflow.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/configure-line-item-workflow.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\igyb53oj.0i3","hash":"/4n/OQoONJzKdwycVjgwEg=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"configure-line-item-workflows\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/organization-administration/configure-line-item-workflow.md\" sourcestartlinenumber=\"26\">Positionsworkflows konfigurieren</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/configure-conditional-decision-workflow.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/configure-conditional-decision-workflow.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\qpexnrwe.txy","hash":"irwZKbf75EUyMZebLJCzBw=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"configure-conditional-decisions-in-a-workflow\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/organization-administration/configure-conditional-decision-workflow.md\" sourcestartlinenumber=\"26\">Konfigurieren von bedingten Entscheidungen in einem Workflow</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/configure-approval-step-workflow.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/configure-approval-step-workflow.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\phng1tws.nyz","hash":"NVbVfc7lUDdyg+qNvx9Bwg=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"configure-approval-steps-in-a-workflow\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/organization-administration/configure-approval-step-workflow.md\" sourcestartlinenumber=\"26\">Genehmigungsschritte in einem Workflow konfigurieren</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/hr/tasks/manage-email-templates.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/hr/tasks/manage-email-templates.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\lv5qccdu.2il","hash":"1THG7AnqNUfslsqZgFIdFQ=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"manage-email-templates\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/hr/tasks/manage-email-templates.md\" sourcestartlinenumber=\"25\">E-Mail-Vorlagen verwalten</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/hr/localizations/tasks/employment-verification-i9-verification.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/hr/localizations/tasks/employment-verification-i9-verification.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\v3u0q4bl.v4k","hash":"5zX+sXq3ZEDDsk1ISFLyGw=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"employment-verification-i9-verification\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/hr/localizations/tasks/employment-verification-i9-verification.md\" sourcestartlinenumber=\"25\">Überprüfung der Beschäftigungsüberprüfung i9</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/saved-views.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/saved-views.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\m5qg5ean.bx5","hash":"AMqChs9ZQ7Zz8eL7TWC/nA=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"saved-views\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/get-started/saved-views.md\" sourcestartlinenumber=\"25\">Gespeicherte Ansichten</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/grid-capabilities.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/grid-capabilities.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\dyqmynm0.bqo","hash":"ugADz2tUeXWmufGjC6w6nA=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"grid-capabilities\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/get-started/grid-capabilities.md\" sourcestartlinenumber=\"25\">Rasterfunktionen</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/client-faq.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/client-faq.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\abh1rms2.jel","hash":"th7SaHC5d7o7MKF/ckEMJg=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"client-faq\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/get-started/client-faq.md\" sourcestartlinenumber=\"26\">Kunden-FAQ</h1>"},{"log_codes":["InvalidFileLink"],"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/MS_Content/index.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/MS_Content/index.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\ksfxnoc0.nbs","hash":"EqzZGKX6CYl1fH0WVp/zjw=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"finance-and-operations-application-documentation\" sourcefile=\"ProcessDoku/00_Basics/MS_Content/index.md\" sourcestartlinenumber=\"26\">Finance and Operations-Anwendungsdokumentation</h1>"},{"log_codes":["InvalidFileLink"],"type":"Conceptual","source_relative_path":"ProcessDoku/00_Basics/Grundlagen_Overview.md","output":{".html":{"relative_path":"ProcessDoku/00_Basics/Grundlagen_Overview.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\z2z4z2s2.upa","hash":"ur0Mfbz4RWRZAQ6zukGYqA=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"benutzeroberfläche-von-d365\" sourcefile=\"ProcessDoku/00_Basics/Grundlagen_Overview.md\" sourcestartlinenumber=\"1\">Benutzeroberfläche von D365</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/03_GlobalDataAndDataExchange/03_02_B2B/B2B_Overview.md","output":{".html":{"relative_path":"ProcessDoku/03_GlobalDataAndDataExchange/03_02_B2B/B2B_Overview.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\fu1ti4ew.jva","hash":"Y8rtm5vdVJJlepW5VGPsMA=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"ProcessDoku/03_GlobalDataAndDataExchange/03_02_B2B/B2B2.md","output":{".html":{"relative_path":"ProcessDoku/03_GlobalDataAndDataExchange/03_02_B2B/B2B2.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\dm4j0kxv.jgx","hash":"1F1zF8Bo+fY6YQfRfQA5TQ=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"ProcessDoku/03_GlobalDataAndDataExchange/03_02_B2B/B2B1.md","output":{".html":{"relative_path":"ProcessDoku/03_GlobalDataAndDataExchange/03_02_B2B/B2B1.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\f5dvzdlx.ps5","hash":"3wJKV/AUtEDqn1HR9+LB9w=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"api/index.md","output":{".html":{"relative_path":"api/index.html","link_to_path":"C:\\D365-Operations\\OwnDocu\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\sd5durkv.hyh","hash":"FTXVsIbwUPdXcrOXXgnFKQ=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"placeholder\" sourcefile=\"api/index.md\" sourcestartlinenumber=\"1\">PLACEHOLDER</h1>"},{"type":"Conceptual","source_relative_path":"index.md","output":{".html":{"relative_path":"index.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\j2baxbas.xlp","hash":"W8kwOKjUCm2sTF0MJHQy4g=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"welcome-to-the-docmentation-of-the-wika-erp-systems-d365\" sourcefile=\"index.md\" sourcestartlinenumber=\"1\">Welcome to the docmentation of the WIKA ERP-Systems D365</h1>"},{"type":"Conceptual","source_relative_path":"ProcessDoku/01_CoreProcesses/01_02_Quotations/Quotations.md","output":{".html":{"relative_path":"ProcessDoku/01_CoreProcesses/01_02_Quotations/Quotations.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\1gnex3sf.he4","hash":"Jy3yxwywoFdPBjvQNe06Nw=="}},"is_incremental":true,"version":"","rawTitle":"<h1 id=\"quotations-overview\" sourcefile=\"ProcessDoku/01_CoreProcesses/01_02_Quotations/Quotations.md\" sourcestartlinenumber=\"5\">Quotations overview</h1>"},{"log_codes":["UidNotFound"],"type":"Conceptual","source_relative_path":"ProcessDoku/01_CoreProcesses/01_03_Sales/Sales_Order.md","output":{".html":{"relative_path":"ProcessDoku/01_CoreProcesses/01_03_Sales/Sales_Order.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\wvxnebyp.1g4","hash":"4pFPBH/+RCCs5mboepbRng=="}},"is_incremental":false,"version":"","rawTitle":"<h1 id=\"create-sales-orders\" sourcefile=\"ProcessDoku/01_CoreProcesses/01_03_Sales/Sales_Order.md\" sourcestartlinenumber=\"5\">Create sales orders</h1>"},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_6.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_6.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_41.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_41.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_3.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_3.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_3.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_29.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_29.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_29.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_51.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_51.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_50.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_50.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_40.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_40.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_4.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_4.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_39.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_39.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_38.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_38.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_31.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_31.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_30.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_30.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/on-hand-inventory.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/on-hand-inventory.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/navigation-search.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/navigation-search.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/lbd-sizing-01.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/lbd-sizing-01.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/keytipsax6.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/keytipsax6.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/howtocontextuallookups-1.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/howtocontextuallookups-1.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/help-pane-ops-help.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/help-pane-ops-help.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/help-architecture.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/help-architecture.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/gridfilteritemlookup.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/gridfilteritemlookup.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/01_03_Sales_Customer_CreateACustTemplate2.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/01_03_Sales_Customer_CreateACustTemplate2.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/01_03_Sales_Customer_CreateACustTemplate2.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/01_03_Sales_Customer_CreateACustTemplate1.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/01_03_Sales_Customer_CreateACustTemplate1.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/01_03_Sales_Customer_CreateACustTemplate1.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/01_03_Sales_Customer_CreateACustTemplate.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/01_03_Sales_Customer_CreateACustTemplate.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/01_03_Sales_Customer_CreateACustTemplate.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/01_03_Sales_Customer_CreateACustomer.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/01_03_Sales_Customer_CreateACustomer.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/01_03_Sales_Customer_CreateACustomer.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/filtereditemlookup.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/filtereditemlookup.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/filtereditemlookup.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/field-description.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/field-description.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/field-description.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_17.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_17.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_16.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_16.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-08.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-08.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-07.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-07.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-02.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-02.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-01.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-01.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/image6.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/image6.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/Create-alert-rule-form.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/Create-alert-rule-form.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/Create-alert-rule-form.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_7.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_7.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/emptyitemlookup.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/emptyitemlookup.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/Create-alert-rule-form.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/Create-alert-rule-form.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/connect-to-lcs-crop.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/connect-to-lcs-crop.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/connect-to-lcs-crop-1024x365.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/connect-to-lcs-crop-1024x365.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/configure-my-workspace.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/configure-my-workspace.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/configure-and-filter-workspaces.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/configure-and-filter-workspaces.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/action-search-field-with-data.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/action-search-field-with-data.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/8c0f12bbb3f26032997ef0ba95d89b6a.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/8c0f12bbb3f26032997ef0ba95d89b6a.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_20.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_20.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_20.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_2.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_2.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_2.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/01_03_Sales_Customer_Texts.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/01_03_Sales_Customer_Texts.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/01_03_Sales_Customer_Texts.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/01_03_Sales_Customer_ExclusiveItem.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/01_03_Sales_Customer_ExclusiveItem.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/01_03_Sales_Customer_ExclusiveItem.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/howtocontextuallookups-1.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/howtocontextuallookups-1.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/howtocontextuallookups-1.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/help-pane-ops-help.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/help-pane-ops-help.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/help-pane-ops-help.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/help-architecture.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/help-architecture.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/help-architecture.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/gridfilteritemlookup.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/gridfilteritemlookup.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/gridfilteritemlookup.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/SalesOrderScheduling.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/SalesOrderScheduling.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/salesandmarketing01.jpg","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/salesandmarketing01.jpg"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/01_03_Sales_Customer_CreateACustTemplate2.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/01_03_Sales_Customer_CreateACustTemplate2.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/01_03_Sales_Customer_CreateACustTemplate1.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/01_03_Sales_Customer_CreateACustTemplate1.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Quotations/NewQuotation_1.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Quotations/NewQuotation_1.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Quotations/NewQuotation.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Quotations/NewQuotation.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Process_Overview_CoreProcesses.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Process_Overview_CoreProcesses.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Process_Map.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Process_Map.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_42.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_42.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_42.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_41.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_41.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_41.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_26.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_26.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_26.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_25.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_25.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_25.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_24.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_24.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_24.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_23.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_23.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_23.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_22.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_22.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_22.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_21.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_21.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_21.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-04.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-04.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-04.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-03.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-03.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-03.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/image4.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/image4.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/image4.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/howtocontextuallookups-2.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/howtocontextuallookups-2.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/howtocontextuallookups-2.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_11.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_11.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_10.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_10.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/01_03_Sales_Customer_CreateACustTemplate.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/01_03_Sales_Customer_CreateACustTemplate.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/01_03_Sales_Customer_CreateACustomer.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/01_03_Sales_Customer_CreateACustomer.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/updatefilterlookupexample.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/updatefilterlookupexample.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/typeaheadlookupexample.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/typeaheadlookupexample.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/rsat-data-agnostic-testing-02.PNG","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/rsat-data-agnostic-testing-02.PNG"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/rsat-data-agnostic-testing-01.PNG","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/rsat-data-agnostic-testing-01.PNG"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/feedback.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/feedback.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/f0d78399e7fafcd85ded1cd1e3d34f3c.jpg","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/f0d78399e7fafcd85ded1cd1e3d34f3c.jpg"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/80f7e8c5ac412fdf2c8a12f7728f135a.jpg","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/80f7e8c5ac412fdf2c8a12f7728f135a.jpg","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/80f7e8c5ac412fdf2c8a12f7728f135a.jpg"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/6d08b0be32808221023e2aa92d69fd70.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/6d08b0be32808221023e2aa92d69fd70.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/6d08b0be32808221023e2aa92d69fd70.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_37.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_37.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_36.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_36.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"images/Production/Ressoucren/00_Ressource_Menu.png","output":{"resource":{"relative_path":"images/Production/Ressoucren/00_Ressource_Menu.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/images/Production/Ressoucren/00_Ressource_Menu.png"}},"is_incremental":false,"version":""},{"type":"Toc","source_relative_path":"toc.yml","output":{".html":{"relative_path":"toc.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\h1dahzfo.zjw","hash":"8zS6TxrZ/Sjbpp3LD9xm9g=="}},"is_incremental":false,"version":""},{"log_codes":["InvalidFileLink"],"type":"Toc","source_relative_path":"api/toc.yml","output":{".html":{"relative_path":"api/toc.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\000p0xik.bye","hash":"OiEFXk7T8Y2AlYcwgbPq6w=="}},"is_incremental":false,"version":""},{"log_codes":["InvalidFileLink"],"type":"Toc","source_relative_path":"ProcessDoku/toc.yml","output":{".html":{"relative_path":"ProcessDoku/toc.html","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365\\obj\\.cache\\build\\2edqtmdf.lnt\\4fexvw4w.505","hash":"nE67HuFPAJYo3LHgzz4RvA=="}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_40.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_40.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_40.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_4.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_4.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_4.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_33.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_33.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_32.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_32.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_28.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_28.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_27.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_27.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_26.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_26.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_25.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_25.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_20.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_20.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_2.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_2.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_19.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_19.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_18.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_18.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/sales01.jpg","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/sales01.jpg"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_34.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_34.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_34.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_19.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_19.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_19.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_18.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_18.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_18.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_17.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_17.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_17.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_16.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_16.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_16.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_15.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_15.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_15.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_14.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_14.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_14.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_13.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_13.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_13.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_12.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_12.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_12.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Quotations/NewQuotation_1.png","output":{"resource":{"relative_path":"ProcessDoku/media/Quotations/NewQuotation_1.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Quotations/NewQuotation_1.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Quotations/NewQuotation.png","output":{"resource":{"relative_path":"ProcessDoku/media/Quotations/NewQuotation.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Quotations/NewQuotation.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Process_Overview_SupportProcesses.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Process_Overview_SupportProcesses.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Process_Overview_GdAndDataExchange.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Process_Overview_GdAndDataExchange.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/organization-administration/media/workflow_multipleusersinstep.gif","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/organization-administration/media/workflow_multipleusersinstep.gif"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/organization-administration/media/workflow_lineitemworkflow.gif","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/organization-administration/media/workflow_lineitemworkflow.gif"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/organization-administration/media/workflow_insertionpoint.gif","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/organization-administration/media/workflow_insertionpoint.gif"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/workspace-section-filters.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/workspace-section-filters.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-06.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-06.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-05.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-05.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-04.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-04.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-03.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-03.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/task-guide-step-1-ops.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/task-guide-step-1-ops.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/task-guide-ops.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/task-guide-ops.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/system-parameters_ops.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/system-parameters_ops.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/system-parameters_ops-1024x437.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/system-parameters_ops-1024x437.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/pages-show-side-by-side.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/pages-show-side-by-side.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/open-in-new-window-icon.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/open-in-new-window-icon.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/media/workflow_insertionpoint.gif","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/media/workflow_insertionpoint.gif","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/organization-administration/media/workflow_insertionpoint.gif"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/workspace-section-filters.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/workspace-section-filters.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/workspace-section-filters.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-02.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-02.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-02.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-01.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-01.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-01.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/updatefilterlookupexample.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/updatefilterlookupexample.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/updatefilterlookupexample.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/typeaheadlookupexample.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/typeaheadlookupexample.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/typeaheadlookupexample.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/pages-show-side-by-side.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/pages-show-side-by-side.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/pages-show-side-by-side.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/open-in-new-window-icon.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/open-in-new-window-icon.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/open-in-new-window-icon.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"images/Prozessübersicht.png","output":{"resource":{"relative_path":"images/Prozessübersicht.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/images/Prozessübersicht.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/images/Picture1.png","output":{"resource":{"relative_path":"docs/images/Picture1.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/marketing01.jpg","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/marketing01.jpg"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/01_03_Sales_Customer_Texts.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/01_03_Sales_Customer_Texts.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/01_03_Sales_Customer_ExclusiveItem.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/01_03_Sales_Customer_ExclusiveItem.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Production/Ressoucren/00_Ressource_Menu.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Production/Ressoucren/00_Ressource_Menu.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Production/Ressoucren/00_Menu_Ressources_gif.gif","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Production/Ressoucren/00_Menu_Ressources_gif.gif"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_28.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_28.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_28.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_27.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_27.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_27.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_11.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_11.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_11.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_10.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_10.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_10.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_1.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_1.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_1.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/SalesOrderScheduling_ReleaseOrder.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/SalesOrderScheduling_ReleaseOrder.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/SalesOrderScheduling_ReleaseOrder.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/SalesOrderScheduling.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/SalesOrderScheduling.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/SalesOrderScheduling.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/salesandmarketing01.jpg","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/salesandmarketing01.jpg","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/salesandmarketing01.jpg"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/sales01.jpg","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/sales01.jpg","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/sales01.jpg"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/marketing01.jpg","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/marketing01.jpg","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/marketing01.jpg"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Basics_Overview.png","output":{"resource":{"relative_path":"ProcessDoku/media/Basics_Overview.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Basics_Overview.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/01_CoreProcesses/01_04_Production/media/ProdPlanningProcess_Overview.png","output":{"resource":{"relative_path":"ProcessDoku/01_CoreProcesses/01_04_Production/media/ProdPlanningProcess_Overview.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/01_CoreProcesses/01_04_Production/media/ProdPlanningProcess_Overview.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/media/workflow_withmanualdecision.gif","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/media/workflow_withmanualdecision.gif","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/organization-administration/media/workflow_withmanualdecision.gif"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/image4.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/image4.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/howtocontextuallookups-2.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/howtocontextuallookups-2.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/filtereditemlookup.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/filtereditemlookup.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/field-description.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/field-description.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/cli-element-property-window.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/cli-element-property-window.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/changingselectionlookup.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/changingselectionlookup.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"images/Picture1.png","output":{"resource":{"relative_path":"images/Picture1.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/images/Picture1.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"images/img1.jpg","output":{"resource":{"relative_path":"images/img1.jpg","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/images/img1.jpg"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/lbd-sizing-01.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/lbd-sizing-01.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/lbd-sizing-01.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/keytipsax6.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/keytipsax6.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/keytipsax6.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"images/Production/Ressoucren/00_Menu_Ressources_gif.gif","output":{"resource":{"relative_path":"images/Production/Ressoucren/00_Menu_Ressources_gif.gif","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/images/Production/Ressoucren/00_Menu_Ressources_gif.gif"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"images/Prozessübersicht AX.png","output":{"resource":{"relative_path":"images/Prozessübersicht AX.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/images/Prozessübersicht AX.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/images/Production/Ressoucren/00_Ressource_Menu.png","output":{"resource":{"relative_path":"docs/images/Production/Ressoucren/00_Ressource_Menu.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/configure-my-workspace.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/configure-my-workspace.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/configure-my-workspace.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/configure-and-filter-workspaces.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/configure-and-filter-workspaces.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/configure-and-filter-workspaces.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/cli-element-property-window.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/cli-element-property-window.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/cli-element-property-window.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/changingselectionlookup.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/changingselectionlookup.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/changingselectionlookup.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/Alert-email-templates.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/Alert-email-templates.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/Alert-email-templates.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/action-search-field.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/action-search-field.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/action-search-field.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_5.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_5.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_49.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_49.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_48.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_48.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_47.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_47.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_46.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_46.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_45.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_45.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_44.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_44.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_43.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_43.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_35.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_35.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_34.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_34.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_5.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_5.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_5.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_49.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_49.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_49.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_33.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_33.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_33.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_32.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_32.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_32.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_31.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_31.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_31.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_30.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_30.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_30.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/image5.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/image5.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/action-search-field-with-data.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/action-search-field-with-data.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/action-search-field-with-data.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/8c0f12bbb3f26032997ef0ba95d89b6a.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/8c0f12bbb3f26032997ef0ba95d89b6a.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/8c0f12bbb3f26032997ef0ba95d89b6a.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_42.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_42.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/personalization-addtoworkspace.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/personalization-addtoworkspace.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/personalization-addtoworkspace.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/connect-to-lcs-crop.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/connect-to-lcs-crop.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/connect-to-lcs-crop.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/connect-to-lcs-crop-1024x365.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/connect-to-lcs-crop-1024x365.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/connect-to-lcs-crop-1024x365.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/fonts/glyphicons-halflings-regular.svg","output":{"resource":{"relative_path":"docs/fonts/glyphicons-halflings-regular.svg"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/logo.svg","output":{"resource":{"relative_path":"docs/logo.svg"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_9.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_9.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_9.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_8.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_8.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_8.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_7.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_7.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_7.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_6.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_6.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_6.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_51.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_51.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_51.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_50.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_50.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_50.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/on-hand-inventory.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/on-hand-inventory.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/on-hand-inventory.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/navigation-search.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/navigation-search.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/navigation-search.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/feedback.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/feedback.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/feedback.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/f0d78399e7fafcd85ded1cd1e3d34f3c.jpg","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/f0d78399e7fafcd85ded1cd1e3d34f3c.jpg","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/f0d78399e7fafcd85ded1cd1e3d34f3c.jpg"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/emptyitemlookup.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/emptyitemlookup.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/emptyitemlookup.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_36.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_36.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_36.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_35.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_35.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_35.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/media/workflow_user.gif","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/media/workflow_user.gif","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/organization-administration/media/workflow_user.gif"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/media/workflow_multipleusersinstep.gif","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/media/workflow_multipleusersinstep.gif","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/organization-administration/media/workflow_multipleusersinstep.gif"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/media/workflow_lineitemworkflow.gif","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/organization-administration/media/workflow_lineitemworkflow.gif","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/organization-administration/media/workflow_lineitemworkflow.gif"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_3.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_3.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_29.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_29.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_24.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_24.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_23.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_23.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_22.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_22.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_21.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_21.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_1.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_1.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/SalesOrderScheduling_ReleaseOrder.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/SalesOrderScheduling_ReleaseOrder.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/images/Prozessübersicht.png","output":{"resource":{"relative_path":"docs/images/Prozessübersicht.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/images/Prozessübersicht AX.png","output":{"resource":{"relative_path":"docs/images/Prozessübersicht AX.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_48.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_48.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_48.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_47.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_47.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_47.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_46.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_46.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_46.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_45.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_45.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_45.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_44.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_44.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_44.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_43.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_43.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_43.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Quotations/Quotation_Scheduling.png","output":{"resource":{"relative_path":"ProcessDoku/media/Quotations/Quotation_Scheduling.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Quotations/Quotation_Scheduling.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Quotations/NewQuotation_2.png","output":{"resource":{"relative_path":"ProcessDoku/media/Quotations/NewQuotation_2.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Quotations/NewQuotation_2.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/workspace-filter.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/workspace-filter.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/workspace-filter.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/workspace-filter-expanded.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/workspace-filter-expanded.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/workspace-filter-expanded.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-08.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-08.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-08.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-07.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-07.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-07.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-06.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-06.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-06.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-05.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-05.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/user-interface-05.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_15.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_15.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_14.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_14.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_13.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_13.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_12.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_12.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Quotations/Quotation_Scheduling.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Quotations/Quotation_Scheduling.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Quotations/NewQuotation_2.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Quotations/NewQuotation_2.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Basics_Overview.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Basics_Overview.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/01_CoreProcesses/01_04_Production/media/ProdPlanningProcess_Overview.png","output":{"resource":{"relative_path":"docs/ProcessDoku/01_CoreProcesses/01_04_Production/media/ProdPlanningProcess_Overview.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/image5.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/image5.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/image5.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/80f7e8c5ac412fdf2c8a12f7728f135a.jpg","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/80f7e8c5ac412fdf2c8a12f7728f135a.jpg"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/images/Production/Ressoucren/00_Menu_Ressources_gif.gif","output":{"resource":{"relative_path":"docs/images/Production/Ressoucren/00_Menu_Ressources_gif.gif"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Production/Ressoucren/00_Ressource_Menu.png","output":{"resource":{"relative_path":"ProcessDoku/media/Production/Ressoucren/00_Ressource_Menu.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Production/Ressoucren/00_Ressource_Menu.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Production/Ressoucren/00_Menu_Ressources_gif.gif","output":{"resource":{"relative_path":"ProcessDoku/media/Production/Ressoucren/00_Menu_Ressources_gif.gif","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Production/Ressoucren/00_Menu_Ressources_gif.gif"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Process_Overview_SupportProcesses.png","output":{"resource":{"relative_path":"ProcessDoku/media/Process_Overview_SupportProcesses.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Process_Overview_SupportProcesses.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Process_Overview_GdAndDataExchange.png","output":{"resource":{"relative_path":"ProcessDoku/media/Process_Overview_GdAndDataExchange.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Process_Overview_GdAndDataExchange.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Process_Overview_CoreProcesses.png","output":{"resource":{"relative_path":"ProcessDoku/media/Process_Overview_CoreProcesses.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Process_Overview_CoreProcesses.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Process_Map.png","output":{"resource":{"relative_path":"ProcessDoku/media/Process_Map.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Process_Map.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/task-guide-step-1-ops.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/task-guide-step-1-ops.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/task-guide-step-1-ops.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/task-guide-ops.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/task-guide-ops.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/task-guide-ops.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/system-parameters_ops.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/system-parameters_ops.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/system-parameters_ops.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/system-parameters_ops-1024x437.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/system-parameters_ops-1024x437.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/system-parameters_ops-1024x437.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/rsat-data-agnostic-testing-02.PNG","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/rsat-data-agnostic-testing-02.PNG","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/rsat-data-agnostic-testing-02.PNG"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/rsat-data-agnostic-testing-01.PNG","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/rsat-data-agnostic-testing-01.PNG","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/rsat-data-agnostic-testing-01.PNG"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/restyledPersonalizationToolbar.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/restyledPersonalizationToolbar.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/restyledPersonalizationToolbar.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/organization-administration/media/workflow_withmanualdecision.gif","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/organization-administration/media/workflow_withmanualdecision.gif"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/organization-administration/media/workflow_user.gif","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/organization-administration/media/workflow_user.gif"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/workspace-filter.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/workspace-filter.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/workspace-filter-expanded.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/workspace-filter-expanded.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/restyledPersonalizationToolbar.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/restyledPersonalizationToolbar.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/personalization-addtoworkspace.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/personalization-addtoworkspace.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/Alert-email-templates.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/Alert-email-templates.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/action-search-field.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/action-search-field.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_9.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_9.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_8.png","output":{"resource":{"relative_path":"docs/ProcessDoku/media/Sales/Guideline/AX2009_8.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/image6.png","output":{"resource":{"relative_path":"ProcessDoku/00_Basics/MS_Content/get-started/media/image6.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/00_Basics/MS_Content/get-started/media/image6.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/6d08b0be32808221023e2aa92d69fd70.png","output":{"resource":{"relative_path":"docs/ProcessDoku/00_Basics/MS_Content/get-started/media/6d08b0be32808221023e2aa92d69fd70.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"docs/images/img1.jpg","output":{"resource":{"relative_path":"docs/images/img1.jpg"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_39.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_39.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_39.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_38.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_38.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_38.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_37.png","output":{"resource":{"relative_path":"ProcessDoku/media/Sales/Guideline/AX2009_37.png","link_to_path":"C:\\Users\\Goldhat\\Documents\\GitHub\\V0_DOKUD365/ProcessDoku/media/Sales/Guideline/AX2009_37.png"}},"is_incremental":false,"version":""}]