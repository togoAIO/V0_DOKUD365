<!DOCTYPE html>
<!--[if IE]><![endif]-->
<html>
  
  <head>
    <meta charset="utf-8">
    <meta http-equiv="X-UA-Compatible" content="IE=edge,chrome=1">
    <title>Configure Accounts receivable and credit and collections | WIKA Documentation </title>
    <meta name="viewport" content="width=device-width">
    <meta name="title" content="Configure Accounts receivable and credit and collections | WIKA Documentation ">
    <meta name="generator" content="docfx 2.56.6.0">
    
    <link rel="shortcut icon" href="../../../../favicon.ico">
    <link rel="stylesheet" href="../../../../styles/docfx.vendor.css">
    <link rel="stylesheet" href="../../../../styles/docfx.css">
    <link rel="stylesheet" href="../../../../styles/main.css">
    <meta property="docfx:navrel" content="../../../../toc.html">
    <meta property="docfx:tocrel" content="../../../toc.html">
    
    <meta property="docfx:rel" content="../../../../">
    
  </head>
  <body data-spy="scroll" data-target="#affix" data-offset="120">
    <div id="wrapper">
      <header>
        
        <nav id="autocollapse" class="navbar navbar-inverse ng-scope" role="navigation">
          <div class="container">
            <div class="navbar-header">
              <button type="button" class="navbar-toggle" data-toggle="collapse" data-target="#navbar">
                <span class="sr-only">Toggle navigation</span>
                <span class="icon-bar"></span>
                <span class="icon-bar"></span>
                <span class="icon-bar"></span>
              </button>
              
              <a class="navbar-brand" href="../../../../index.html">
                <img id="logo" class="svg" src="../../../../logo.svg" alt="">
              </a>
            </div>
            <div class="collapse navbar-collapse" id="navbar">
              <form class="navbar-form navbar-right" role="search" id="search">
                <div class="form-group">
                  <input type="text" class="form-control" id="search-query" placeholder="Search" autocomplete="off">
                </div>
              </form>
            </div>
          </div>
        </nav>
        
        <div class="subnav navbar navbar-default">
          <div class="container hide-when-search" id="breadcrumb">
            <ul class="breadcrumb">
              <li></li>
            </ul>
          </div>
        </div>
      </header>
      <div class="container body-content">
        
        <div id="search-results">
          <div class="search-list">Search Results for <span></span></div>
          <div class="sr-items">
            <p><i class="glyphicon glyphicon-refresh index-loading"></i></p>
          </div>
          <ul id="pagination" data-first="First" data-prev="Previous" data-next="Next" data-last="Last"></ul>
        </div>
      </div>
      <div role="main" class="container body-content hide-when-search">
        
        <div class="sidenav hide-when-search">
          <a class="btn toc-toggle collapse" data-toggle="collapse" href="#sidetoggle" aria-expanded="false" aria-controls="sidetoggle">Show / Hide Table of Contents</a>
          <div class="sidetoggle collapse" id="sidetoggle">
            <div id="sidetoc"></div>
          </div>
        </div>
        <div class="article row grid-right">
          <div class="col-md-10">
            <article class="content wrap" id="_content" data-uid="">
<h1 id="configure-accounts-receivable-and-credit-and-collections" sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="30">Configure Accounts receivable and credit and collections</h1>

[!include[banner](../includes/banner.md)]
<p sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="34">Configure Accounts receivable and Credit and Collections to track invoices and incoming payments from customers.</p>
<p sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="36">You can set up customer groups, customers, posting profiles, various payment options, interest notes, collection letters, commissions, parameters regarding customers, charges, deliveries and destinations, bills of exchange, and other types of Accounts receivable and Credit and collections information.
The following table lists the pages that support the configuration and maintenance of Accounts receivable and Credit and collections. The table entries are organized by task and then alphabetically by page name.</p>
<div class="NOTE" sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="39">
<h5>Note</h5>
<p sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="40">You cannot navigate to some pages in the following table unless data or parameter settings have been entered in other pages.</p>
</div>
<table sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="42">
<thead>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="42">
<th sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="42">Task</th>
<th sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="42">Page name</th>
<th sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="42">Usage</th>
</tr>
</thead>
<tbody>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="44">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="44">Configuring required Accounts receivable information</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="44">Accounts receivable parameters</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="44">Set up parameters for the Accounts receivable module.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="45">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="45"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="45">Accounts receivable workflows</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="45">Create a workflow or modify an existing one.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="46">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="46"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="46">Customer groups</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="46">Create and maintain groups of customers who share key parameters. These include terms of payment, settle periods, inventory posting ledger accounts, sales tax group, and default account setup.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="47">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="47"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="47">Customer posting profile</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="47">Set up the posting profiles that control the posting of customer transactions to the general ledger.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="48">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="48"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="48">Form setup</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="48">Define the format of information on various documents that are related to customers, such as sales orders, picking lists, packing slips, and invoices.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="49">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="49"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="49">Methods of payment - customer</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="49">Create and maintain information about methods of payment for customers.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="50">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="50"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="50">Terms of payment</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="50">Define the terms of payment that you assign to sales orders, purchase orders, customers, and vendors in either Accounts receivable or Accounts payable.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="51">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="51"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="51"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="51"></td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="52">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="52">Configuring Accounts receivable journals</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="52">Journal names</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="52">Create and manage templates for journals. This includes the management of posting restrictions for selected users or user groups.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="53">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="53"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="53"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="53"></td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="54">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="54">Configuring customer invoices</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="54">Billing codes</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="54">Set up optional codes for billing charges to use on free text invoice lines.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="55">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="55"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="55">Charges code</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="55">Set up codes for the charges to use on sales orders and purchase orders, such as invoice fees, freight, and insurance.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="56">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="56"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="56">Footer text</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="56">Specify footer text for a print management record in multiple languages. When the document is printed, the language of the document determines the language of the footer text.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="57">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="57"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="57">Form notes</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="57">Edit the standard text that appears on the various pages that your organization uses, such as invoices, sales orders, and interest notes.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="58">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="58"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="58">Form setup</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="58">Define page note parameters for quotations, confirmations, picking lists, packing slips, customer invoices, free text invoices, and interest notes.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="59">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="59"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="59">Form sorting parameters</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="59">Set up sorting orders for printing multiple invoices, such as by invoice account and sales order number.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="60">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="60"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="60">Print management setup</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="60">Set up print management original or copy records and conditional settings. This information controls the way that documents, such as sales orders and purchase orders, are printed during the confirmation process.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="61">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="61"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="61"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="61"></td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="62">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="62">Configuring customer payments</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="62">Cash discounts</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="62">Set up and manage cash discount codes, which are linked to customer and vendor accounts and are applied to sales orders and purchase orders.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="63">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="63"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="63">Credit card processors</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="63">Set up information for credit card processors that authorize credit cards that are submitted for the payment of sales orders.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="64">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="64"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="64">Currencies</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="64">Create and view the currencies that your organization uses.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="65">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="65"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="65">Currency exchange rates</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="65">Create and maintain appropriate exchange rates between the accounting currency and other currencies.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="66">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="66"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="66">Intercompany accounting</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="66">Create a list of accounts that the current legal entity can post to. You must set up debit and credit accounts, and also set up the journal that receives the transactions in the other legal entity.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="67">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="67"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="67">Methods of payment - customer</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="67">Create and maintain information about methods of payment for customers. For more information, see <a href="tasks/establish-customer-method-payment.html" sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="67">Establish customer method of payment</a>.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="68">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="68"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="68">Organization hierarchies</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="68">Set up an organization hierarchy for centralized payments.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="69">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="69"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="69">Organization hierarchy purposes</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="69">Specify a purpose for centralized payments.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="70">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="70"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="70">Payment days</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="70">Define the payment days that are used to calculate due dates for payments that you will receive from customers or make to vendors.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="71">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="71"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="71">Payment fee</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="71">Create and maintain payment fees that are related to customers, such as fees for bills of exchange.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="72">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="72"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="72">Payment fee setup</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="72">Set up payment fees for various combinations of banks, methods of payment, remittance types, payment specifications, currencies, and date intervals.  For more information, see <a href="tasks/establish-customer-payment-fees.html" sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="72">Establish customer payment fees</a>.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="73">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="73"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="73">Payment schedules</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="73">Create payment schedules, which you can use to schedule installment payments from customers and to vendors.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="74">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="74"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="74">Payment specification</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="74">Create and view payment specification codes for the method of payment that you selected in the Methods of payment page. You define payment specification codes according to your agreement with the bank that is specified for the selected method of payment.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="75">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="75"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="75">Transaction text</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="75">Create transaction text for automatic postings to General ledger. You can set up transaction text in various languages.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="76">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="76"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="76">Translations</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="76">Create text in another language. You can translate all texts for external use (such as terms of payment, terms of delivery, and modes of delivery) into one or more languages.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="77">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="77"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="77"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="77"></td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="78">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="78">Configuring customer payment formats</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="78">Bill of exchange layout</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="78">Set up the layout of bills of exchange for the bank account that you selected in the Bank accounts page.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="79">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="79"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="79">Check layout</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="79">Set up the layout of checks for the bank account that you selected in the Bank accounts page.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="80">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="80"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="80">File formats for methods of payment</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="80">Select import, export, return, and remittance file formats to use for customer payments.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="81">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="81"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="81">Methods of payment - customer</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="81">Create and maintain information about methods of payment for customers.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="82">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="82"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="82">Signature</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="82">Add, change, or remove signature image files, such as .bmp, .jpg, or .gif files. The signature image files are printed on checks as official legal entity signatures.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="83">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="83"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="83"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="83"></td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="84">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="84">Configuring Accounts receivable statistics</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="84">Aging period definitions</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="84">Set up and manage user-defined aging period definitions, which are used to analyze the maturity of customer accounts and vendor accounts, based on a date that you enter. For more information, see <a href="tasks/set-up-accounts-receivable-aging-information.html" sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="84">Set up and generate accounts receivable aging information</a>.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="85">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="85"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="85">Business statistics</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="85">Set up business statistics inquiries that can help you analyze the performance of your organization.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="86">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="86"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="86">Business statistics data</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="86">View data in a grid format for a selected business statistic.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="87">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="87"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="87"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="87"></td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="88">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="88">Maintaining customer information</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="88">Address book</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="88">Enter or view information about prospects, leads, opportunities, customers, contact persons, competitors, and employees.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="89">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="89"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="89">Customer bank accounts</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="89">Create and manage customer bank accounts.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="90">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="90"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="90">Customer groups</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="90">Create and maintain groups of customers who share key parameters. These include terms of payment, settle periods, inventory posting ledger accounts, sales tax group, and default account setup.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="91">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="91"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="91">Customers</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="91">Create and manage the customer accounts for the customers the organization does business with.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="92">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="92"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="92">Print management setup</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="92">Set up print management original or copy records and conditional settings. This information controls the way that documents, such as sales orders and purchase orders, are printed during the posting process.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="93">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="93"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="93"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="93"></td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="94">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="94">Configuring Credit and collections</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="94">Accounts receivable parameters</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="94">Set up parameters for the Credit and Collections module.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="95">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="95"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="95">Case categories</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="95">Set up a case category that will be used for Collections cases.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="96">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="96"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="96">Collection letter</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="96">Create and manage collection letter sequences and connect them with collection letter lines.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="97">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="97"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="97">Collections agent</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="97">Set up collections agents for use in the Collections page.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="98">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="98"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="98">Collections team</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="98">Set up a collections team that represents the workers that can be setup as agents. A team called Collections will be setup automatically in the Accounts receivable parameters if no team exists.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="99">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="99"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="99">Customer aging snapshot</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="99">Create aging snapshots for customers. An aging snapshot contains the calculated aged balances for a group of customers at one point in time. This step requires an aging period definition to be setup.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="100">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="100"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="100">Customer contacts and email settings</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="100">Set up contacts for customers with their email addresses. These addresses will appear in the Collections page and will be used to create emails that go to customers. Also set up a default Collections contact for each customer that will appear first in the Collections page.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="101">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="101"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="101">Customer pools</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="101">Set up customer pools, which are queries that define a group of customer accounts that can be displayed and managed for collections or aging processes.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="102">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="102"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="102">Customer posting profile</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="102">Set up the profiles that control the posting of customer transactions to the general ledger.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="103">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="103"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="103">Customer reason codes</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="103">Set up customer reasons codes.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="104">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="104"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="104">Customer write-off reason codes</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="104">Set up customer write-off reasons codes that will be used for write-off transactions.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="105">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="105"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="105">Form setup</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="105">Define form note parameters for quotations, confirmations, picking lists, packing slips, customer invoices, free text invoices, and interest notes.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="106">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="106"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="106">Interest</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="106">Set up and manage interest codes.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="107">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="107"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="107">NSF information.</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="107">Set up NSF information on the bank account that will be used when a payment is marked as an NSF transaction on the Collections page.</td>
</tr>
<tr sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="108">
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="108"></td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="108">Salesperson information</td>
<td sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="108">Set up the email address for salespersons. These addresses will appear on the Collections page and you can use them to send email to a salesperson from that page.</td>
</tr>
</tbody>
</table>
<p sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="111">For more information, see <a href="collections-credit-accounts-receivable.html" sourcefile="ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md" sourcestartlinenumber="111">Credit and collections in Accounts receivable</a>.</p>
[!include[footer-include](../../includes/footer-banner.md)]</article>
          </div>
          
          <div class="hidden-sm col-md-2" role="complementary">
            <div class="sideaffix">
              <div class="contribution">
                <ul class="nav">
                  <li>
                    <a href="https://github.com/togoAIO/V0_DOKUD365/blob/master/ProcessDoku/02_SupportProcesses/02_01_Finance/accounts-receivable/accounts-receivables-set-up-overview.md/#L1" class="contribution-link">Improve this Doc</a>
                  </li>
                </ul>
              </div>
              <nav class="bs-docs-sidebar hidden-print hidden-xs hidden-sm affix" id="affix">
                <h5>In This Article</h5>
                <div></div>
              </nav>
            </div>
          </div>
        </div>
      </div>
      
      <footer>
        <div class="grad-bottom"></div>
        <div class="footer">
          <div class="container">
            <span class="pull-right">
              <a href="#top">Back to top</a>
            </span>
            <span>Customized Footer</span>
            
          </div>
        </div>
      </footer>
    </div>
    
    <script type="text/javascript" src="../../../../styles/docfx.vendor.js"></script>
    <script type="text/javascript" src="../../../../styles/docfx.js"></script>
    <script type="text/javascript" src="../../../../styles/main.js"></script>
  </body>
</html>
