a   �
  a   v   ]  z  a  n  �  �  e  z  �  �  �     	   	  ,	  :	  F	  b	  �
  �
     v   FileAndType�   ]  �{"baseDir":"C:/Users/Goldhat/Documents/GitHub/V0_DOKUD365","file":"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md","type":"article","sourceDir":"","destinationDir":""}   z  OriginalFileAndType�   a  �{"baseDir":"C:/Users/Goldhat/Documents/GitHub/V0_DOKUD365","file":"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md","type":"article","sourceDir":"","destinationDir":""}   n  Keyo   �  e~/ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md   �  LocalPathFromRootm   e  cProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md   z  LinkToFiles   �  �  �  d  g   �  ]~/ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites.mdn   d  d~/ProcessDoku/02_SupportProcesses/fin-ops-core/dev-itpro/data-entities/configure-export-data-lake.mdf   �  \~/ProcessDoku/02_SupportProcesses/fin-ops-core/fin-ops/imp-lifecycle/environment-planning.md   �  
LinkToUids	   �        FileLinkSources  	  �{"~/ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites.md":[{"Target":"~/ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites.md","SourceFile":"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md","LineNumber":38}],"~/ProcessDoku/02_SupportProcesses/fin-ops-core/dev-itpro/data-entities/configure-export-data-lake.md":[{"Target":"~/ProcessDoku/02_SupportProcesses/fin-ops-core/dev-itpro/data-entities/configure-export-data-lake.md","SourceFile":"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md","LineNumber":69}],"~/ProcessDoku/02_SupportProcesses/fin-ops-core/fin-ops/imp-lifecycle/environment-planning.md":[{"Target":"~/ProcessDoku/02_SupportProcesses/fin-ops-core/fin-ops/imp-lifecycle/environment-planning.md","SourceFile":"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md","LineNumber":45}]}    	  UidLinkSources   ,	  {}   :	  Uids   F	  []   b	  ManifestPropertiesm  �
  �{"rawTitle":"<h1 id=\"configuration-for-finance-insights-for-public-preview-preview---version-10020-and-later\" sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"29\">Configuration for Finance insights for public preview (preview) - version 10.0.20 and later</h1>"}   �
  DocumentType	   �
   �� o� {"$type":"System.Collections.Generic.Dictionary`2[[System.String, mscorlib],[System.Object, mscorlib]], mscorlib","conceptual":"\n[!include[rename-banner](~/includes/cc-data-platform-banner.md)]\n<p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"35\">Finance insights combines functionality from Microsoft Dynamics 365 Finance with Dataverse, Azure, and AI Builder to provide powerful forecasting tools for your organization. This topic explains how to configure Dynamics 365 Finance version 10.0.20 so that your system can use the capabilities that are available in Finance insights public preview.</p>\n<div class=\"NOTE\" sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"37\">\n<h5>Note</h5>\n<p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"38\">The configuration steps that are described in this topic apply only to Finance version 10.0.20 and later. 'To set up Finance insights on version 10.0.19 and earlier, see <a href=\"~/ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites.md\" sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"38\">Configuration for Finance insights - versions up to 10.0.19</a>.</p>\n</div>\n<h2 id=\"deploy-finance\" sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"40\">Deploy Finance</h2>\n<p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"42\">Follow these steps to deploy the environments.</p>\n<ol sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"44\">\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"44\">In Microsoft Dynamics Lifecycle Services (LCS), create or update a Finance environment. The environment requires app version 10.0.20 or later of Finance and Operations apps.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"45\">The environment must be a high-availability (HA) environment in Sandbox. (This type of environment is also known as a Tier-2 environment.) For more information, see <a href=\"../../fin-ops-core/fin-ops/imp-lifecycle/environment-planning.md\" sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"45\">Environment planning</a>.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"46\">If you are configuring Finance insights in a Sandbox environment, you might need to copy production data to that environment for predictions to work. The prediction model uses multiple years of data to build predictions. The Contoso demo data doesn’t contain enough historical data to train the prediction model adequately.</li>\n</ol>\n<h2 id=\"configure-dataverse\" sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"48\">Configure Dataverse</h2>\n<p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"50\">Follow these steps to configure Dataverse for Finance insights.</p>\n<ol sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"52\">\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"52\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"52\">In LCS, open the environment page, and verify that the <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"52\">Power Platform Integration</strong> section is already set up.</p>\n<ul sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"54\">\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"54\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"54\">If it's already set up, the Dataverse environment name that is linked to the Finance environment should be listed.</p>\n</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"55\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"55\">If it isn't yet set up, follow these steps:</p>\n<ol sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"57\">\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"57\">In the <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"57\">Power Platform Integration</strong> section, select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"57\">Setup</strong>. Setup of the environment might take up to an hour.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"58\">If the Dataverse environment is successfully set up, the Dataverse environment name that is linked to the Finance environment should be listed.</li>\n</ol>\n<div class=\"NOTE\" sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"60\">\n<h5>Note</h5>\n<p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"61\">After you complete the environment setup, do <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"61\">not</strong> select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"61\">Link to CDS for Apps</strong>. This button isn't required for Finance insights. If you select it, you won't be able to configure the required environment add-ins in LCS.</p>\n</div>\n</li>\n</ul>\n</li>\n</ol>\n<h2 id=\"configure-azure\" sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"63\">Configure Azure</h2>\n<h3 id=\"use-azure-cloud-shell-to-set-up-finance-insights-data-lake-resources\" sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"65\">Use Azure Cloud Shell to set up Finance insights Data Lake resources</h3>\n<div class=\"tabGroup\" id=\"tabgroup_CeZOj-G++Q\" sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"67\">\n<ul role=\"tablist\">\n<li role=\"presentation\">\n<a href=\"#tabpanel_CeZOj-G++Q_use-a-powershell-script\" role=\"tab\" aria-controls=\"tabpanel_CeZOj-G++Q_use-a-powershell-script\" data-tab=\"use-a-powershell-script\" tabindex=\"0\" aria-selected=\"true\" sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"67\">Use a Windows PowerShell script</a>\n</li>\n<li role=\"presentation\">\n<a href=\"#tabpanel_CeZOj-G++Q_azure-azure-cli\" role=\"tab\" aria-controls=\"tabpanel_CeZOj-G++Q_azure-azure-cli\" data-tab=\"azure-azure-cli\" tabindex=\"-1\" sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"222\">Azure CLI</a>\n</li>\n</ul>\n<section id=\"tabpanel_CeZOj-G++Q_use-a-powershell-script\" role=\"tabpanel\" data-tab=\"use-a-powershell-script\">\n\n<p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"69\">A Windows PowerShell script has been provided so that you can easily set up the Azure resources that are described in <a href=\"../../fin-ops-core/dev-itpro/data-entities/configure-export-data-lake.md\" sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"69\">Configure export to Azure Data Lake</a>. If you prefer to do the setup manually, skip this procedure, and complete the procedure in the <a href=\"#manual-setup\" sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"69\">Manual setup</a> section instead.</p>\n<div class=\"NOTE\" sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"71\">\n<h5>Note</h5>\n<p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"72\">Use the following procedure to run the Windows PowerShell script. The setup might not work if you use the <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"72\">Try it</strong> option in Azure CLI or if you run the script on your computer.</p>\n</div>\n<p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"74\">Follow these steps to use the Windows PowerShell script to configure Azure. You must have rights to create an Azure resource group, Azure resources, and an Azure AD application. For information about the required permissions, see <a href=\"/azure/active-directory/develop/howto-create-service-principal-portal#permissions-required-for-registering-an-app\" sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"74\">Check Azure AD permissions</a>.</p>\n<ol sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"76\">\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"76\">In the <a href=\"https://portal.azure.com\" sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"76\">Azure portal</a>, go to your target Azure subscription.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"77\">Select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"77\">Cloud Shell</strong> to the right of the <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"77\">Search</strong> field.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"78\">Select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"78\">PowerShell</strong>.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"79\">Create storage if you're prompted to create it.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"80\">On the <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"80\">Azure CLI</strong> tab, select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"80\">Copy</strong>.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"81\">In Notepad, open a new file, and paste in the Windows PowerShell script.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"82\">Save the file as <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"82\">ConfigureDataLake.ps1</strong>.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"83\">Upload the Windows PowerShell script to the session by using the menu option for upload in Cloud Shell.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"84\">Run the <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"84\">.\\ConfigureDataLake.ps1</strong> script.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"85\">Follow the prompts to run the script.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"86\">Use the information from the script output to install the Export to Data Lake add-in in LCS.</li>\n</ol>\n<h3 id=\"manual-setup\" sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"88\">Manual setup</h3>\n<h4 id=\"add-applications-to-the-azure-ad-tenant\" sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"90\">Add applications to the Azure AD tenant</h4>\n<ol sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"92\">\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"92\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"92\">In the <a href=\"https://portal.azure.com\" sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"92\">Azure portal</a>, go to <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"92\">Azure Active Directory</strong>.</p>\n</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"93\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"93\">Select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"93\">Manage &gt; Enterprise applications</strong>.</p>\n</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"94\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"94\">Search for the following applications by app ID.</p>\n<table sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"96\">\n<thead>\n<tr sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"96\">\n<th sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"96\">Application</th>\n<th sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"96\">App ID</th>\n</tr>\n</thead>\n<tbody>\n<tr sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"98\">\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"98\">Microsoft Dynamics ERP Microservices</td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"98\">0cdb527f-a8d1-4bf8-9436-b352c68682b2</td>\n</tr>\n<tr sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"99\">\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"99\">Microsoft Dynamics ERP Microservices CDS</td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"99\">703e2651-d3fc-48f5-942c-74274233dba8</td>\n</tr>\n<tr sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"100\">\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"100\">AI Builder Authorization Service</td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"100\">ad40333e-9910-4b61-b281-e3aeeb8c3ef3</td>\n</tr>\n</tbody>\n</table>\n</li>\n</ol>\n<p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"102\">If you can't find any of the preceding applications, try the following steps.</p>\n<ol sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"104\">\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"104\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"104\">On your local computer, on the <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"104\">Start</strong> menu, search for <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"104\">powershell</strong>.</p>\n</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"105\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"105\">Select and hold (or right-click) <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"105\">Windows PowerShell</strong>, and then select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"105\">Run as administrator</strong>.</p>\n</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"106\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"106\">Run the following command to install the <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"106\">AzureAD</strong> module.</p>\n<p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"108\"><code sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"108\">Install-Module -Name AzureAD</code></p>\n</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"110\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"110\">If a NuGet provider is required to continue, select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"110\">Y</strong> to install it.</p>\n</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"111\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"111\">If you receive an &quot;Untrusted repository&quot; message, select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"111\">Y</strong> to continue.</p>\n</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"112\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"112\">For each application that must be added, run the following commands to add the application to Azure AD. When you're prompted, sign in as the Azure AD administrator.</p>\n<p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"114\"><code sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"114\">Connect-AzureAD</code></p>\n<p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"116\"><code sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"116\">New-AzureADServicePrincipal –AppId &lt;AppId&gt;</code></p>\n</li>\n</ol>\n<h4 id=\"create-azure-resources\" sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"118\">Create Azure resources</h4>\n<div class=\"NOTE\" sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"120\">\n<h5>Note</h5>\n<p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"121\">Make sure that you create the following resources in the same Azure AD instance that the Dataverse environment is in. You can't use resources from a different Azure AD instance.</p>\n</div>\n<ol sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"123\">\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"123\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"123\">Create a storage account:</p>\n<ol sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"125\">\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"125\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"125\">In the <a href=\"https://portal.azure.com\" sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"125\">Azure portal</a>, create a storage account.</p>\n</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"126\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"126\">In the <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"126\">Create storage account</strong> dialog box, set the following fields:</p>\n<ul sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"128\">\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"128\"><strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"128\">Location</strong> – Select the data center where your environment is located.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"129\"><strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"129\">Performance</strong> – We recommend that you select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"129\">Standard</strong>.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"130\"><strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"130\">Account kind</strong> – You must select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"130\">StorageV2</strong>.</li>\n</ul>\n</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"132\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"132\">In the <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"132\">Advanced options</strong> dialog box, for the <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"132\">Data Lake storage Gen2</strong> option, select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"132\">Enable</strong> under the <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"132\">Hierarchical namespaces</strong> feature. If you don't enable this feature, you can't consume data that Finance and Operations apps write by using services such as Power BI data flows.</p>\n</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"133\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"133\">Select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"133\">Review and create</strong>. When the deployment is completed, the new resource is shown in the Azure portal.</p>\n</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"134\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"134\">Go to the storage account that you created.</p>\n</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"135\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"135\">On the left menu, select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"135\">Access keys</strong>.</p>\n</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"136\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"136\">Copy and save the name of the storage account. You will have to provide this value later, when you set up key vault secrets.</p>\n</li>\n</ol>\n</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"138\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"138\">Create a key vault:</p>\n<ol sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"140\">\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"140\">In the <a href=\"https://portal.azure.com\" sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"140\">Azure portal</a>, create a key vault.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"141\">In the <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"141\">Create key vault</strong> dialog box, in the <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"141\">Location</strong> field, select the data center where your environment is located.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"142\">After key vault is created, go to <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"142\">Key Vault Overview</strong>, and copy and save the DNS name. You will have to provide this value later, when you set up the Data Lake add-in.</li>\n</ol>\n</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"144\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"144\">Create and register an Azure AD application:</p>\n<ol sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"146\">\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"146\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"146\">In the <a href=\"https://portal.azure.com\" sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"146\">Azure portal</a>, go to <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"146\">Azure Active Directory</strong>, and then select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"146\">App registrations</strong>.</p>\n</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"147\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"147\">Select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"147\">New application registration</strong>, and set the following fields:</p>\n<ul sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"149\">\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"149\"><strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"149\">Name</strong> – Enter the name of the app.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"150\"><strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"150\">Application type</strong> – Select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"150\">Web API</strong>.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"151\"><strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"151\">Redirect URI setup</strong> – Enter the URL for your Dynamics 365 instance, such as <code sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"151\">https://yourdynamicsinstance.dynamics.com/auth</code>.</li>\n</ul>\n</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"153\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"153\">Go to the app that you just created, and copy and save its <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"153\">Application (client) ID</strong> value. You will have to provide this value later, when you set up key vault secrets.</p>\n</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"154\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"154\">Go to <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"154\">API permissions</strong>, and follow these steps:</p>\n<ol sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"156\">\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"156\">Select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"156\">Add a permission</strong>.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"157\">Select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"157\">Azure Key vault</strong>.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"158\">After you select delegated permissions, select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"158\">user_impersonation</strong>.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"159\">Select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"159\">Add permissions</strong>.</li>\n</ol>\n</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"161\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"161\">On the menu for the app, select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"161\">Certificates &amp; secrets</strong>, and then follow these steps to create Key Vault secrets:</p>\n<ol sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"163\">\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"163\">Select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"163\">New client secret</strong>.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"164\">In the <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"164\">Key Description</strong> field, enter a name.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"165\">Select a duration, and then select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"165\">Add</strong>. A secret is generated in the <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"165\">Value</strong> field.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"166\">Copy and save the client secret value. You will have to provide this value later, when you set up key vault secrets.</li>\n</ol>\n</li>\n</ol>\n</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"168\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"168\">Create Key Vault secrets:</p>\n<ol sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"170\">\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"170\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"170\">Go to the key vault that you created earlier, and select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"170\">Secrets</strong>.</p>\n</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"171\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"171\">For each secret name in the following table, follow these steps:</p>\n<ol sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"173\">\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"173\">Select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"173\">Generate/Import</strong>.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"174\">In the <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"174\">Create a secret</strong> dialog box, in the <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"174\">Upload options</strong> field, select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"174\">Manual</strong>.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"175\">Create the secret name and value from the table.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"176\">Select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"176\">Enabled</strong>, and then select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"176\">Create</strong>. The secret is created and added to Key Vault.</li>\n</ol>\n<table sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"178\">\n<thead>\n<tr sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"178\">\n<th sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"178\">Secret name</th>\n<th sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"178\">Secret value</th>\n</tr>\n</thead>\n<tbody>\n<tr sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"180\">\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"180\">app-id</td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"180\">The app ID of the application that you created earlier.</td>\n</tr>\n<tr sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"181\">\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"181\">app-secret</td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"181\">The client secret that you saved earlier.</td>\n</tr>\n<tr sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"182\">\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"182\">storage-account-name</td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"182\">The name of the storage account that you created earlier, such as <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"182\">storageaccount1</strong>.</td>\n</tr>\n</tbody>\n</table>\n</li>\n</ol>\n</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"184\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"184\">Authorize the application to access the key vault:</p>\n<ol sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"186\">\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"186\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"186\">In the <a href=\"https://portal.azure.com\" sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"186\">Azure portal</a>, open the key vault that you created earlier.</p>\n</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"187\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"187\">Select the access policies.</p>\n</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"188\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"188\">For each application in the following table, follow these steps:</p>\n<ol sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"190\">\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"190\">Select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"190\">Add Access Policy</strong> to create an access policy.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"191\">In the <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"191\">Secret permissions</strong> field, select the permissions from the table.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"192\">In the <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"192\">Select principal</strong> field, search for the application display name from the table.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"193\">Select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"193\">Select</strong>.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"194\">Select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"194\">Add</strong>.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"195\">Select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"195\">Save</strong>.</li>\n</ol>\n<table sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"197\">\n<thead>\n<tr sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"197\">\n<th sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"197\">Application</th>\n<th sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"197\">Permissions</th>\n</tr>\n</thead>\n<tbody>\n<tr sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"199\">\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"199\">The display name of the new application that you created</td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"199\">Get, List</td>\n</tr>\n<tr sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"200\">\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"200\"><strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"200\">Microsoft Dynamics ERP Microservices</strong></td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"200\">Get, List</td>\n</tr>\n</tbody>\n</table>\n</li>\n</ol>\n</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"202\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"202\">Assign roles to access the storage account:</p>\n<ol sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"204\">\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"204\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"204\">In the <a href=\"https://portal.azure.com\" sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"204\">Azure portal</a>, open the storage account that you created earlier.</p>\n</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"205\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"205\">Select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"205\">Access Control (IAM)</strong>, and then select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"205\">Role Assignments</strong>.</p>\n</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"206\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"206\">Select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"206\">Add, Add Role Assignment</strong>.</p>\n</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"207\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"207\">For each application in the following table, follow these steps:</p>\n<ol sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"209\">\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"209\">Select the role from the table.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"210\">Leave the <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"210\">Assign access to</strong> field set to <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"210\">Azure AD user, group, or service principal</strong>.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"211\">In the <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"211\">Select</strong> field, enter the application from the table.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"212\">Select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"212\">Save</strong>.</li>\n</ol>\n<table sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"214\">\n<thead>\n<tr sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"214\">\n<th sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"214\">Application</th>\n<th sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"214\">Role</th>\n</tr>\n</thead>\n<tbody>\n<tr sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"216\">\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"216\">The display name of the new application that you created</td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"216\">Owner</td>\n</tr>\n<tr sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"217\">\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"217\">The display name of the new application that you created</td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"217\">Contributor</td>\n</tr>\n<tr sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"218\">\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"218\">The display name of the new application that you created</td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"218\">Storage Account Contributor</td>\n</tr>\n<tr sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"219\">\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"219\">The display name of the new application that you created</td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"219\">Storage Blob Data Owner</td>\n</tr>\n<tr sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"220\">\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"220\"><strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"220\">AI Builder Authorization Service</strong></td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"220\">Storage Blob Data Reader</td>\n</tr>\n</tbody>\n</table>\n</li>\n</ol>\n</li>\n</ol>\n</section>\n<section id=\"tabpanel_CeZOj-G++Q_azure-azure-cli\" role=\"tabpanel\" data-tab=\"azure-azure-cli\" aria-hidden=\"true\" hidden=\"hidden\">\n\n<pre><code sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"224\">function New-FinanceDataLakeAzureResources {\n    Assert-ScriptSetup\n\n    $ClientAppName = 'Finance Data Lake Application'\n    $DefaultSecretExpiryInYear = 1\n    $MicrosoftDynamicsERPMicroservicesAppId = '0cdb527f-a8d1-4bf8-9436-b352c68682b2'\n    $MicrosoftDynamicsERPMicroservicesCDSAppId = '703e2651-d3fc-48f5-942c-74274233dba8'\n    $AIBuilderAuthorizationServiceAppId = 'ad40333e-9910-4b61-b281-e3aeeb8c3ef3'\n    $KeyVaultServicePrincipalAppId = 'cfa8b339-82a2-471a-a3c9-0fc0be7a4093'\n    $GraphServicePrincipalAppId = '00000003-0000-0000-c000-000000000000'\n\n    Import-Module AzureAD.Standard.Preview\n    $connectAzureADParameters = @{ 'Identity' = $true; 'TenantId' = $env:ACC_TID }\n    $azContext = AzureAD.Standard.Preview\\Connect-AzureAD @connectAzureADParameters\n    $userContext = ConvertFrom-Json ((az ad signed-in-user show) -join '')\n    $user = Get-AzureADUser -Filter (&quot;UserPrincipalName eq '&quot; + $userContext.UserPrincipalName + &quot;'&quot;)\n\n    Set-AzureSubscription\n    \n    $resourceGroup = $null\n    $ResourceGroupName = 'D365FinanceInsightsDataLake'\n    $ResourceGroupNameSuffix = ''\n    $FullResourceGroupName = ''\n    Write-Output (&quot;The default Azure Resource Group name is '{0}'&quot; -f $ResourceGroupName)\n    while (-not ($resourceGroup)) {\n        $ResourceGroupNameSuffix = (Read-Host -Prompt &quot;Enter optional Azure Resource Group name suffix: (leave blank for no suffix)&quot;)\n        if ([string]::IsNullOrWhitespace($ResourceGroupNameSuffix))\n        {\n            $FullResourceGroupName = $ResourceGroupName\n        }\n        else\n        {\n            if ($ResourceGroupNameSuffix -notmatch &quot;^[A-Za-z0-9]+$&quot;) {\n                Write-Warning &quot;The Azure Resource Group name suffix can only include alphanumeric characters.&quot;\n                continue\n            }\n\n            if ($ResourceGroupNameSuffix.Length -gt 60) {\n                Write-Warning &quot;The Azure Resource Group name suffix cannot be longer than 60 characters.&quot;\n                continue\n            }\n\n            $FullResourceGroupName = $ResourceGroupName + $ResourceGroupNameSuffix\n        }\n        \n        $resourceGroup = Get-AzResourceGroup -Name $FullResourceGroupName -ErrorAction SilentlyContinue\n\n        if (-not ($resourceGroup)) {\n            Write-Output (&quot;Your new Azure Resource Group name is '{0}'&quot; -f $FullResourceGroupName)\n            $resourceLocation = ''\n            $azResourceLocations = (Get-AzLocation | Select-Object Location).Location\n            while ([string]::IsNullOrWhitespace($resourceLocation) -or (-not ($resourceLocation -in $azResourceLocations))) {\n                $resourceLocation = (Read-Host -Prompt &quot;Enter the location in which to create the Azure Resource Group: ('help' to see values)&quot;)\n                if ($resourceLocation -eq 'help') {\n                    Write-Output (&quot;List of available regions is '{0}'&quot; -f ($azResourceLocations -join ','))\n                }\n                elseif ([string]::IsNullOrWhitespace($resourceLocation) -or (-not ($resourceLocation -in $azResourceLocations)))\n                {\n                    Write-Warning (&quot;The provided location is not available for resource group. List of available regions is '{0}'&quot; -f ($azResourceLocations -join ','))\n                }\n            }\n            $resourceGroup = New-AzResourceGroup -Name $FullResourceGroupName -Location $resourceLocation\n            Write-Output (&quot;Created Azure Resource Group '{0}'&quot; -f $resourceGroup.ResourceGroupName)\n        }\n        else {\n            Write-Output (&quot;Found Azure Resource Group '{0}'&quot; -f ($resourceGroup.ResourceGroupName))\n        }\n    }\n\n    Write-Output '================================================================================='\n    $MicrosoftDynamicsERPMicroservicesAppObjectId = Create-ADServicePrincipal -AppId $MicrosoftDynamicsERPMicroservicesAppId\n    Create-ADServicePrincipal -AppId $MicrosoftDynamicsERPMicroservicesCDSAppId | Out-Null\n    $aibuilderAuthorizationServiceObjectId = Create-ADServicePrincipal -AppId $AIBuilderAuthorizationServiceAppId\n    Write-Output ('=================================================================================')\n\n    $clientAppSPN = Get-AzureADServicePrincipal -Filter (&quot;DisplayName eq '&quot; + $ClientAppName + &quot;'&quot;)\n    if (-not ($clientAppSPN)) {\n        $keyVaultPrincipal = Get-AzureADServicePrincipal -Filter (&quot;AppId eq '&quot; + $KeyVaultServicePrincipalAppId + &quot;'&quot;)\n        if (-not $keyVaultPrincipal)\n        {\n            New-AzureADServicePrincipal -AppId $KeyVaultServicePrincipalAppId | Format-Table -AutoSize\n            Write-Output &quot;Added Key Vault principal to AAD&quot;\n            $keyVaultPrincipal = Get-AzureADServicePrincipal -Filter (&quot;AppId eq '&quot; + $KeyVaultServicePrincipalAppId + &quot;'&quot;)\n        }\n        $keyVaultAccess = New-Object -TypeName &quot;Microsoft.Open.AzureAD.Model.RequiredResourceAccess&quot;\n        $keyVaultAccess.ResourceAppId = $keyVaultPrincipal.AppId\n        $keyVaultAccess.ResourceAccess = (New-Object -TypeName &quot;microsoft.open.azuread.model.resourceAccess&quot; -ArgumentList $keyVaultPrincipal.Oauth2Permissions.Id, &quot;Scope&quot;)\n\n        $graphPrincipal = Get-AzureADServicePrincipal -Filter (&quot;AppId eq '&quot; + $GraphServicePrincipalAppId + &quot;'&quot;)\n        if (-not $graphPrincipal)\n        {\n            New-AzureADServicePrincipal -AppId $GraphServicePrincipalAppId | Format-Table -AutoSize\n            Write-Output &quot;Added Graph principal to AAD&quot;\n            $graphPrincipal = Get-AzureADServicePrincipal -Filter (&quot;AppId eq '&quot; + $GraphServicePrincipalAppId + &quot;'&quot;)\n        }\n        $userRead = $graphPrincipal.Oauth2Permissions | Where-Object { $_.Type -eq &quot;User&quot; -and $_.Value -eq &quot;User.Read&quot; }\n        $graphAccess = New-Object -TypeName &quot;Microsoft.Open.AzureAD.Model.RequiredResourceAccess&quot;\n        $graphAccess.ResourceAppId = $graphPrincipal.AppId\n        $graphAccess.ResourceAccess = (New-Object -TypeName &quot;microsoft.open.azuread.model.resourceAccess&quot; -ArgumentList $userRead.Id, &quot;Scope&quot;)\n\n        $clientApp = New-AzureADApplication -DisplayName $ClientAppName -RequiredResourceAccess @($keyVaultAccess, $graphAccess)\n        $clientAppSPN = New-AzureADServicePrincipal -AppId $clientApp.AppId -Tags @($ClientAppName)\n        $clientAppId = $clientApp.AppId\n        Write-Output ('Created App Registration &quot;' + $ClientAppName + '&quot; with Application Id: ' + $clientAppId)\n    }\n    else {\n        $clientApp = Get-AzureADApplication -Filter (&quot;DisplayName eq '&quot; + $ClientAppName + &quot;'&quot;)\n        $clientAppId = $clientApp.AppId\n        Write-Output ('Found App Registration &quot;' + $ClientAppName + '&quot; with Application Id: ' + $clientAppId)\n    }\n            \n    $clientAppSecretCredential = New-AzureADApplicationPasswordCredential -ObjectId $clientApp.ObjectId -CustomKeyIdentifier &quot;ClientAppAccessKey&quot; -EndDate (get-date).AddYears($DefaultSecretExpiryInYear)\n    $ClientAppSecret = $clientAppSecretCredential.Value\n    $clientAppSpId = $clientAppSPN.ObjectId\n\n    Write-Output ('Generated application secret: ' + $ClientAppSecret)\n    Write-Output '================================================================================='\n\n    $templateObject = ConvertFrom-Json $azureTemplate -AsHashtable\n    $templateObject.{$schema} = &quot;https://schema.management.azure.com/schemas/2019-04-01/deploymentTemplate.json#&quot;\n    Write-Output 'Provisioning Azure resources. This may take a few minutes.'\n    try {\n        $deployment = New-AzResourceGroupDeployment -ResourceGroupName $FullResourceGroupName -TemplateObject $templateObject -aibuilderAppObjectId $aibuilderAuthorizationServiceObjectId -clientAppId $clientAppId -clientAppSecret $ClientAppSecret -clientAppSpObjectId  $clientAppSpId -microserviceSpObjectId $MicrosoftDynamicsERPMicroservicesAppObjectId -userSpObjectId $user.ObjectId -Force -ErrorAction Stop\n    }\n    catch {\n        $ErrorMessage = $_.Exception.Message\n        if ($ErrorMessage.Contains(&quot;not allowed to be updated&quot;))\n        {\n            Write-Error ($ErrorMessage)\n            Write-Warning &quot;Some items in the existing resource group $FullResourceGroupName could not be updated. To resolve the issue, remove the existing resource group $FullResourceGroupName and run the script again.&quot;\n        }\n        else {\n            throw\n        }\n\n    }\n    if ($deployment.ProvisioningState -eq 'Succeeded') {\n        Write-Output &quot;Successfully deployed the following resources to Azure:&quot;\n        Write-Output (&quot;  Key Vault:                         &quot; + $deployment.Outputs.keyVaultName.Value)\n        Write-Output (&quot;  Storage Account:                   &quot; + $deployment.Outputs.storageAccountName.Value)\n        \n        $keyVault = Get-AzKeyVault -VaultName $deployment.Outputs.keyVaultName.Value\n        $tenantId = (Get-AzContext).Tenant.Id\n\n        Write-Output &quot;Values for LCS Data Lake Add-In:&quot;\n        Write-Output (&quot;  Tenant ID:                         &quot; + $tenantId)\n        Write-Output (&quot;  DNS Name:                          &quot; + $keyVault.VaultUri)\n        Write-Output &quot;  Storage account secret name:       storage-account-name&quot;\n        Write-Output &quot;  Application ID secret name:        app-id&quot;\n        Write-Output &quot;  Application Secret secret name:    app-secret&quot;\n        Write-Warning &quot;Copy this information for the LCS Add-in for easy access. Azure Cloud Shell will eventually time out and close.&quot;\n\n        Write-Output '================================================================================='\n        Write-Output &quot;Values for System parameters &gt; Data connections:&quot;\n        Write-Output (&quot;  Application ID:                    &quot; + $clientAppId)\n        Write-Output (&quot;  Application Secret:                &quot; + $ClientAppSecret)\n        Write-Output (&quot;  DNS name:                          &quot; + $keyVault.VaultUri)\n        Write-Output &quot;  Secret name:                       storage-account-connection-string&quot;\n        Write-Warning &quot;Copy this information for the System parameters for easy access. Azure Cloud Shell will eventually time out and close.&quot;\n    }\n    else {\n        Write-Output (&quot;Provisioning Azure resources failed with the following state: &quot; + $deployment.ProvisioningState)\n        Write-Output (&quot;Some of the resources may have been created in resource group: &quot; + $FullResourceGroupName)\n    }\n}\n\nfunction Assert-ScriptSetup {\n    if ($PSVersionTable.PSEdition -ne 'Core' -or -not $env:ACC_TID) { \n        throw &quot;This script needs to be uploaded and run from Azure Cloud Shell (PowerShell).&quot; \n    }\n    \n    if ((Get-AzContext) -eq $null -and (Connect-AzAccount) -eq $null) {\n        throw 'Unable to connect to Azure account.'\n    }\n}\n\nfunction Set-AzureSubscription {\n    $azSubscription = $null\n    while (-not ($azSubscription)) {\n        $subscriptionId = (Read-Host -Prompt &quot;Enter the Azure Subscription ID: (leave blank for default)&quot;)\n        if ([string]::IsNullOrWhitespace($subscriptionId)){\n            break\n        }\n        elseif (-not [guid]::TryParse($subscriptionId, $([ref][guid]::Empty))) {\n                Write-Warning &quot;Azure Subscription ID must be a valid GUID.&quot;\n                continue\n        }\n\n        $azSubscription = Select-AzSubscription -SubscriptionId $subscriptionId\n    }\n}\n\nfunction Create-ADServicePrincipal {\n    param (\n        [string] $AppId\n    )\n\n    $service = Get-AzureADServicePrincipal -Filter (&quot;AppId eq '&quot; + $AppId + &quot;'&quot;)\n    if (-not $service) {\n        New-AzureADServicePrincipal -AppId $AppId | Out-Null\n        $service = Get-AzureADServicePrincipal -Filter (&quot;AppId eq '&quot; + $AppId + &quot;'&quot;)\n        Write-Host (&quot;Added AAD Enterprise Application {0} with Application ID {1}&quot; -f $service.DisplayName,$AppId)\n    }\n    else {\n        Write-Host (&quot;Found AAD Enterprise Application {0} with Application ID {1}&quot; -f $service.DisplayName,$AppId)\n    }\n\n    return $service.ObjectId\n}\n\n$azureTemplate = @&quot;\n{\n    &quot;contentVersion&quot;: &quot;1.0.0.0&quot;,\n    &quot;parameters&quot;: {\n      &quot;aibuilderAppObjectId&quot;: {\n        &quot;type&quot;: &quot;string&quot;,\n        &quot;metadata&quot;: {\n          &quot;description&quot;: &quot;Specifies the object ID of the AI Builder application.&quot;\n        }\n      },\n      &quot;clientAppId&quot;: {\n        &quot;type&quot;: &quot;string&quot;,\n        &quot;metadata&quot;: {\n          &quot;description&quot;: &quot;Specifies the application ID of client application.&quot;\n        }\n      },\n      &quot;clientAppSecret&quot;: {\n        &quot;type&quot;: &quot;String&quot;,\n        &quot;metadata&quot;: {\n          &quot;description&quot;: &quot;Specifies the Azure App ID client secret to in azure key vault.&quot;\n        }\n      },\n      &quot;clientAppSpObjectId&quot;: {\n        &quot;type&quot;: &quot;string&quot;,\n        &quot;metadata&quot;: {\n          &quot;description&quot;: &quot;Specifies the object ID of a client application service principal.&quot;\n        }\n      },\n      &quot;userSpObjectId&quot;: {\n        &quot;type&quot;: &quot;string&quot;,\n        &quot;metadata&quot;: {\n          &quot;description&quot;: &quot;Specifies the object ID of tenant admin service principal.&quot;\n        }\n      },\n      &quot;microserviceSpObjectId&quot;: {\n        &quot;type&quot;: &quot;string&quot;,\n        &quot;metadata&quot;: {\n          &quot;description&quot;: &quot;Specifies the object ID of Microsoft Dynamics ERP Microservices service principal.&quot;\n        }\n      },\n      &quot;storageAccountType&quot;: {\n        &quot;type&quot;: &quot;string&quot;,\n        &quot;defaultValue&quot;: &quot;Standard_LRS&quot;,\n        &quot;allowedValues&quot;: [\n          &quot;Standard_LRS&quot;,\n          &quot;Standard_GRS&quot;,\n          &quot;Standard_ZRS&quot;,\n          &quot;Premium_LRS&quot;\n        ],\n        &quot;metadata&quot;: {\n          &quot;description&quot;: &quot;Storage Account type&quot;\n        }\n      }\n    },\n    &quot;variables&quot;: {\n      &quot;storageAccountApiVersion&quot;: &quot;2019-06-01&quot;,\n      &quot;keyVaultApiVersion&quot;: &quot;2018-02-14&quot;,\n      &quot;secretsPermissions&quot;: [\n        &quot;list&quot;,\n        &quot;get&quot;\n      ],\n      &quot;location&quot;: &quot;[resourceGroup().location]&quot;,\n      &quot;storageAccountName&quot;: &quot;[concat('store', uniquestring(resourceGroup().id))]&quot;,\n      &quot;keyVaultName&quot;: &quot;[concat('keyvault', uniquestring(resourceGroup().id))]&quot;,\n      &quot;owner&quot;: &quot;[concat('/subscriptions/', subscription().subscriptionId, '/providers/Microsoft.Authorization/roleDefinitions/', '8e3af657-a8ff-443c-a75c-2fe8c4bcb635')]&quot;,\n      &quot;contributor&quot;: &quot;[concat('/subscriptions/', subscription().subscriptionId, '/providers/Microsoft.Authorization/roleDefinitions/', 'b24988ac-6180-42a0-ab88-20f7382dd24c')]&quot;,\n      &quot;storageAccountContributor&quot;: &quot;[concat('/subscriptions/', subscription().subscriptionId, '/providers/Microsoft.Authorization/roleDefinitions/', '17d1049b-9a84-46fb-8f53-869881c3d3ab')]&quot;,\n      &quot;storageBlobDataOwner&quot;: &quot;[concat('/subscriptions/', subscription().subscriptionId, '/providers/Microsoft.Authorization/roleDefinitions/', 'b7e6dc6d-f1e8-4753-8033-0f276bb0955b')]&quot;,\n      &quot;storageBlobDataReader&quot;: &quot;[concat('/subscriptions/', subscription().subscriptionId, '/providers/Microsoft.Authorization/roleDefinitions/', '2a2b9908-6ea1-4ae2-8e65-a410df84e7d1')]&quot;\n    },\n    &quot;resources&quot;: [\n      {\n        &quot;type&quot;: &quot;Microsoft.Storage/storageAccounts&quot;,\n        &quot;apiVersion&quot;: &quot;[variables('storageAccountApiVersion')]&quot;,\n        &quot;name&quot;: &quot;[variables('storageAccountName')]&quot;,\n        &quot;location&quot;: &quot;[variables('location')]&quot;,\n        &quot;sku&quot;: {\n          &quot;name&quot;: &quot;[parameters('storageAccountType')]&quot;\n        },\n        &quot;kind&quot;: &quot;StorageV2&quot;,\n        &quot;properties&quot;: {\n          &quot;accessTier&quot;: &quot;Hot&quot;,\n          &quot;supportsHttpsTrafficOnly&quot;: true,\n          &quot;isHnsEnabled&quot;: true\n        },\n        &quot;resources&quot;: [\n          {\n            &quot;type&quot;: &quot;Microsoft.Storage/storageAccounts/providers/roleAssignments&quot;,\n            &quot;apiVersion&quot;: &quot;2018-09-01-preview&quot;,\n            &quot;name&quot;: &quot;[concat(variables('storageAccountName'), '/Microsoft.Authorization/', guid(uniqueString(variables('storageAccountName'),'1')))]&quot;,\n            &quot;dependsOn&quot;: [\n              &quot;[variables('storageAccountName')]&quot;\n            ],\n            &quot;properties&quot;: {\n              &quot;roleDefinitionId&quot;: &quot;[variables('owner')]&quot;,\n              &quot;principalId&quot;: &quot;[parameters('clientAppSpObjectId')]&quot;\n            }\n          },\n          {\n            &quot;type&quot;: &quot;Microsoft.Storage/storageAccounts/providers/roleAssignments&quot;,\n            &quot;apiVersion&quot;: &quot;2018-09-01-preview&quot;,\n            &quot;name&quot;: &quot;[concat(variables('storageAccountName'), '/Microsoft.Authorization/', guid(uniqueString(variables('storageAccountName'),'2')))]&quot;,\n            &quot;dependsOn&quot;: [\n              &quot;[variables('storageAccountName')]&quot;\n            ],\n            &quot;properties&quot;: {\n              &quot;roleDefinitionId&quot;: &quot;[variables('contributor')]&quot;,\n              &quot;principalId&quot;: &quot;[parameters('clientAppSpObjectId')]&quot;\n            }\n          },\n          {\n            &quot;type&quot;: &quot;Microsoft.Storage/storageAccounts/providers/roleAssignments&quot;,\n            &quot;apiVersion&quot;: &quot;2018-09-01-preview&quot;,\n            &quot;name&quot;: &quot;[concat(variables('storageAccountName'), '/Microsoft.Authorization/', guid(uniqueString(variables('storageAccountName'),'3')))]&quot;,\n            &quot;dependsOn&quot;: [\n              &quot;[variables('storageAccountName')]&quot;\n            ],\n            &quot;properties&quot;: {\n              &quot;roleDefinitionId&quot;: &quot;[variables('storageAccountContributor')]&quot;,\n              &quot;principalId&quot;: &quot;[parameters('clientAppSpObjectId')]&quot;\n            }\n          },\n          {\n            &quot;type&quot;: &quot;Microsoft.Storage/storageAccounts/providers/roleAssignments&quot;,\n            &quot;apiVersion&quot;: &quot;2018-09-01-preview&quot;,\n            &quot;name&quot;: &quot;[concat(variables('storageAccountName'), '/Microsoft.Authorization/', guid(uniqueString(variables('storageAccountName'),'4')))]&quot;,\n            &quot;dependsOn&quot;: [\n              &quot;[variables('storageAccountName')]&quot;\n            ],\n            &quot;properties&quot;: {\n              &quot;roleDefinitionId&quot;: &quot;[variables('storageBlobDataOwner')]&quot;,\n              &quot;principalId&quot;: &quot;[parameters('clientAppSpObjectId')]&quot;\n            }\n          },\n          {\n            &quot;type&quot;: &quot;Microsoft.Storage/storageAccounts/providers/roleAssignments&quot;,\n            &quot;apiVersion&quot;: &quot;2018-09-01-preview&quot;,\n            &quot;name&quot;: &quot;[concat(variables('storageAccountName'), '/Microsoft.Authorization/', guid(uniqueString(variables('storageAccountName'),'5')))]&quot;,\n            &quot;dependsOn&quot;: [\n              &quot;[variables('storageAccountName')]&quot;\n            ],\n            &quot;properties&quot;: {\n              &quot;roleDefinitionId&quot;: &quot;[variables('storageBlobDataReader')]&quot;,\n              &quot;principalId&quot;: &quot;[parameters('aibuilderAppObjectId')]&quot;\n            }\n          }\n        ]\n      },\n      {\n        &quot;type&quot;: &quot;Microsoft.KeyVault/vaults&quot;,\n        &quot;apiVersion&quot;: &quot;[variables('keyVaultApiVersion')]&quot;,\n        &quot;name&quot;: &quot;[variables('keyVaultName')]&quot;,\n        &quot;location&quot;: &quot;[variables('location')]&quot;,\n        &quot;dependsOn&quot;: [\n          &quot;[resourceId('Microsoft.Storage/storageAccounts', variables('storageAccountName'))]&quot;\n        ],\n        &quot;tags&quot;: {\n        },\n        &quot;properties&quot;: {\n          &quot;enabledForDeployment&quot;: false,\n          &quot;enabledForTemplateDeployment&quot;: false,\n          &quot;enabledForDiskEncryption&quot;: false,\n          &quot;enableRbacAuthorization&quot;: false,\n          &quot;accessPolicies&quot;: [\n            {\n              &quot;objectId&quot;: &quot;[parameters('clientAppSpObjectId')]&quot;,\n              &quot;tenantId&quot;: &quot;[subscription().tenantId]&quot;,\n              &quot;permissions&quot;: {\n                &quot;secrets&quot;: &quot;[variables('secretsPermissions')]&quot;\n              }\n            },\n            {\n              &quot;objectId&quot;: &quot;[parameters('microserviceSpObjectId')]&quot;,\n              &quot;tenantId&quot;: &quot;[subscription().tenantId]&quot;,\n              &quot;permissions&quot;: {\n                &quot;secrets&quot;: &quot;[variables('secretsPermissions')]&quot;\n              }\n            },\n            {\n              &quot;objectId&quot;: &quot;[parameters('userSpObjectId')]&quot;,\n              &quot;tenantId&quot;: &quot;[subscription().tenantId]&quot;,\n              &quot;permissions&quot;: {\n                &quot;secrets&quot;: &quot;[variables('secretsPermissions')]&quot;\n              }\n            }\n          ],\n          &quot;tenantId&quot;: &quot;[subscription().tenantId]&quot;,\n          &quot;sku&quot;: {\n            &quot;name&quot;: &quot;Standard&quot;,\n            &quot;family&quot;: &quot;A&quot;\n          },\n          &quot;enableSoftDelete&quot;: false,\n          &quot;networkAcls&quot;: {\n            &quot;defaultAction&quot;: &quot;Allow&quot;,\n            &quot;bypass&quot;: &quot;AzureServices&quot;\n          }\n        }\n      },\n      {\n        &quot;type&quot;: &quot;Microsoft.KeyVault/vaults/secrets&quot;,\n        &quot;name&quot;: &quot;[concat(variables('keyVaultName'), '/', 'app-id')]&quot;,\n        &quot;apiVersion&quot;: &quot;[variables('keyVaultApiVersion')]&quot;,\n        &quot;location&quot;: &quot;[variables('location')]&quot;,\n        &quot;dependsOn&quot;: [\n          &quot;[resourceId('Microsoft.KeyVault/vaults', variables('keyVaultName'))]&quot;\n        ],\n        &quot;properties&quot;: {\n          &quot;value&quot;: &quot;[parameters('clientAppId')]&quot;\n        }\n      },\n      {\n        &quot;type&quot;: &quot;Microsoft.KeyVault/vaults/secrets&quot;,\n        &quot;name&quot;: &quot;[concat(variables('keyVaultName'), '/', 'app-secret')]&quot;,\n        &quot;apiVersion&quot;: &quot;[variables('keyVaultApiVersion')]&quot;,\n        &quot;location&quot;: &quot;[variables('location')]&quot;,\n        &quot;dependsOn&quot;: [\n          &quot;[resourceId('Microsoft.KeyVault/vaults', variables('keyVaultName'))]&quot;\n        ],\n        &quot;properties&quot;: {\n          &quot;value&quot;: &quot;[parameters('clientAppSecret')]&quot;\n        }\n      },\n      {\n        &quot;type&quot;: &quot;Microsoft.KeyVault/vaults/secrets&quot;,\n        &quot;name&quot;: &quot;[concat(variables('keyVaultName'), '/', 'storage-account-name')]&quot;,\n        &quot;apiVersion&quot;: &quot;[variables('keyVaultApiVersion')]&quot;,\n        &quot;location&quot;: &quot;[variables('location')]&quot;,\n        &quot;dependsOn&quot;: [\n          &quot;[resourceId('Microsoft.KeyVault/vaults', variables('keyVaultName'))]&quot;\n        ],\n        &quot;properties&quot;: {\n          &quot;value&quot;: &quot;[variables('storageAccountName')]&quot;\n        }\n      },\n      {\n        &quot;type&quot;: &quot;Microsoft.KeyVault/vaults/secrets&quot;,\n        &quot;name&quot;: &quot;[concat(variables('keyVaultName'), '/', 'storage-account-connection-string')]&quot;,\n        &quot;apiVersion&quot;: &quot;[variables('keyVaultApiVersion')]&quot;,\n        &quot;location&quot;: &quot;[variables('location')]&quot;,\n        &quot;dependsOn&quot;: [\n          &quot;[resourceId('Microsoft.KeyVault/vaults', variables('keyVaultName'))]&quot;\n        ],\n        &quot;properties&quot;: {\n          &quot;value&quot;: &quot;[concat('DefaultEndpointsProtocol=https;AccountName=', variables('storageAccountName'), ';AccountKey=', listKeys(resourceId('Microsoft.Storage/storageAccounts', variables('storageAccountName')), variables('storageAccountApiVersion')).keys[0].value, ';EndpointSuffix=core.windows.net')]&quot;\n        }\n      }\n    ],\n    &quot;outputs&quot;: {\n      &quot;storageAccountName&quot;: {\n        &quot;type&quot;: &quot;string&quot;,\n        &quot;value&quot;: &quot;[variables('storageAccountName')]&quot;\n      },\n      &quot;keyVaultName&quot;: {\n        &quot;type&quot;: &quot;string&quot;,\n        &quot;value&quot;: &quot;[variables('keyVaultName')]&quot;\n      }\n    }\n  }\n&quot;@\n\ntry {\n  Start-Transcript -path (Join-Path $HOME Provision-FinInsights-Azure.log)\n  New-FinanceDataLakeAzureResources\n}\ncatch {\n  Write-Error $_.Exception.Message\n\n  if ($PSItem.Exception.StackTrace -ne $null)\n  {\n      Write-Warning $_.Exception.StackTrace\n  }\n\n  $inner = $_.Exception.InnerException\n  while ($null -ne $inner) {\n    Write-Output 'Inner Exception:'\n    Write-Error $_.Exception.Message\n    Write-Warning $_.Exception.StackTrace\n    $inner = $inner.InnerException\n  }\n}\nfinally {\n  Stop-Transcript\n}\n</code></pre>\n</section>\n</div>\n<h2 id=\"configure-the-export-to-data-lake-add-in\" sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"721\">Configure the Export to Data Lake add-in</h2>\n<p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"723\">Follow these steps to use LCS to add the Export to Data Lake add-in to the environment.</p>\n<ol sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"725\">\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"725\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"725\">Sign in to LCS, and then, under the environment name on the right side of the page, select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"725\">Full Details</strong>.</p>\n</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"726\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"726\">In the <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"726\">Environment add-ins</strong> section, select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"726\">Install a new add-in</strong>.</p>\n</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"727\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"727\">Select the <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"727\">Export to Data Lake</strong> add-in.</p>\n</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"728\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"728\">Enter the following values.</p>\n<table sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"730\">\n<thead>\n<tr sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"730\">\n<th sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"730\">Value</th>\n<th sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"730\">Description</th>\n</tr>\n</thead>\n<tbody>\n<tr sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"732\">\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"732\">Tenant ID of the Azure Subscription where the Key Vault is located</td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"732\">The tenant ID where the storage account, apps, and key vaults are located. To obtain this value, open the <a href=\"https://portal.azure.com\" sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"732\">Azure portal</a>, go to <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"732\">Azure Active Directory</strong>, and copy the <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"732\">Tenant ID</strong> value.</td>\n</tr>\n<tr sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"733\">\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"733\">Provide the DNS name of your Key Vault</td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"733\">The DNS name of the key vault, such as <code sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"733\">https://customkeyvault.vault.azure.net/</code>.</td>\n</tr>\n<tr sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"734\">\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"734\">Provide the secret that contains the name of the storage account</td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"734\"><strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"734\">storage-account-name</strong></td>\n</tr>\n<tr sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"735\">\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"735\">Secret Name for App ID to be used for accessing Data Lake</td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"735\"><strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"735\">app-id</strong></td>\n</tr>\n<tr sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"736\">\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"736\">Secret name for App client secret</td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"736\"><strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"736\">app-secret</strong></td>\n</tr>\n</tbody>\n</table>\n</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"738\"><p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"738\">Agree to the terms, and then select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"738\">Install</strong>.</p>\n</li>\n</ol>\n<p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"740\">The add-in will be installed within a few minutes.</p>\n<h2 id=\"configure-the-finance-insights-add-in\" sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"742\">Configure the Finance insights add-in</h2>\n<div class=\"NOTE\" sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"744\">\n<h5>Note</h5>\n<p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"745\">If you previously installed the Get insights add-in, uninstall it before you complete the following procedure.</p>\n</div>\n<p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"747\">Follow these steps to install the Finance insights add-in.</p>\n<ol sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"749\">\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"749\">Sign in to LCS, and then, under the environment name on the right side of the page, select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"749\">Full Details</strong>.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"750\">In the <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"750\">Environment add-ins</strong> section, select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"750\">Install a new add-in</strong>.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"751\">Select the <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"751\">Finance insights</strong> add-in.</li>\n<li sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"752\">Agree to the terms, and then select <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"752\">Install</strong>.</li>\n</ol>\n<p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"754\">The add-in might take several minutes to install.</p>\n<h2 id=\"feedback-and-support\" sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"756\">Feedback and support</h2>\n<p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"758\">If you're interested in providing feedback, or if you require support, send an email to <a href=\"mailto:fiap@microsoft.com\" sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"758\">Finance insights (Preview)</a>.</p>\n[!include[footer-include](../../includes/footer-banner.md)]","type":"Conceptual","source":{"$type":"Microsoft.DocAsCode.DataContracts.Common.SourceDetail, Microsoft.DocAsCode.DataContracts.Common","remote":{"$type":"Microsoft.DocAsCode.Common.Git.GitDetail, Microsoft.DocAsCode.Common","path":"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md","branch":"master","repo":"https://github.com/togoAIO/V0_DOKUD365.git"},"startLine":0,"endLine":0,"isExternal":false},"path":"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md","documentation":{"$type":"Microsoft.DocAsCode.DataContracts.Common.SourceDetail, Microsoft.DocAsCode.DataContracts.Common","remote":{"$type":"Microsoft.DocAsCode.Common.Git.GitDetail, Microsoft.DocAsCode.Common","path":"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md","branch":"master","repo":"https://github.com/togoAIO/V0_DOKUD365.git"},"startLine":0,"endLine":0,"isExternal":false},"_enableSearch":"true","_docfxVersion":"2.56.6.0","_appTitle":"WIKA Documentation","_systemKeys":{"$type":"System.String[], mscorlib","$values":["conceptual","type","source","path","documentation","title","rawTitle","wordCount"]},"rawTitle":"<h1 id=\"configuration-for-finance-insights-for-public-preview-preview---version-10020-and-later\" sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/finance-insights/configure-for-fin-insites-PubPrvw.md\" sourcestartlinenumber=\"29\">Configuration for Finance insights for public preview (preview) - version 10.0.20 and later</h1>","ms.custom":14151,"title":"Configuration for Finance insights for public preview (preview) - version 10.0.20 and later","ms.dyn365.ops.version":"AX 10.0.20","ms.search.region":"Global","ms.assetid":"3d43ba40-780c-459a-a66f-9a01d556e674","author":"ShivamPandey-msft","description":"This topic explains how to configure your system to use the capabilities that are available in Finance insights for public preview in version 10.0.20 and later.","ms.author":"shpandey","audience":"Application User","ms.search.validFrom":"2021-06-03","ms.topic":"article","ms.search.form":null,"ms.date":"06/16/2021","ms.technology":null,"ms.prod":null,"ms.reviewer":"roschlom"}�   � {"$type":"System.Collections.Generic.Dictionary`2[[System.String, mscorlib],[System.Object, mscorlib]], mscorlib","IsUserDefinedTitle":true,"XrefSpec":null}	   �  