a   )  a   v   ]  z  a  n  �  �  e  z  �  �  �  �  �  �  �  �      
        v   FileAndType�   ]  �{"baseDir":"C:/Users/Goldhat/Documents/GitHub/V0_DOKUD365","file":"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md","type":"article","sourceDir":"","destinationDir":""}   z  OriginalFileAndType�   a  �{"baseDir":"C:/Users/Goldhat/Documents/GitHub/V0_DOKUD365","file":"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md","type":"article","sourceDir":"","destinationDir":""}   n  Keyo   �  e~/ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md   �  LocalPathFromRootm   e  cProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md   z  LinkToFiles	   �     �  
LinkToUids	   �     �  FileLinkSources   �  {}   �  UidLinkSources   �  {}   �  Uids     []     ManifestProperties�   
  �{"rawTitle":"<h1 id=\"standard-payroll-reports\" sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"30\">Standard payroll reports</h1>"}      DocumentType	   )   >  9C  {"$type":"System.Collections.Generic.Dictionary`2[[System.String, mscorlib],[System.Object, mscorlib]], mscorlib","conceptual":"\n[!include[banner](../../includes/banner.md)]\n<p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"34\">This topic describes the standard payroll reports that are provided to help you with payroll processing and government reporting. Use these standard reports to create pay statements and W-2 forms that you can issue to your workers, validate payroll taxes and benefit amounts, and complete federal and state regulatory reports.</p>\n<p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"36\">This topic describes functionality that is available only if the <strong sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"36\">Payroll - USA</strong> configuration key is selected.</p>\n<h2 id=\"payroll-standard-reports\" sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"38\">Payroll standard reports</h2>\n<p sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"40\">The following table summarizes when and why you use each report.</p>\n<table sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"42\">\n<thead>\n<tr sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"42\">\n<th sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"42\">Report</th>\n<th sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"42\">Every pay period</th>\n<th sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"42\">Quarterly</th>\n<th sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"42\">Annually</th>\n<th sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"42\">As required</th>\n</tr>\n</thead>\n<tbody>\n<tr sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"44\">\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"44\">Pay statements</td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"44\">After you generate the payroll payment journal, use this report to print pay statements that you can issue to workers.</td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"44\"></td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"44\"></td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"44\">Use this report to reprint pay statements for workers.</td>\n</tr>\n<tr sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"45\">\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"45\">Benefit register</td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"45\">Use this report to validate the benefit amounts that were calculated during payroll processing.</td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"45\"></td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"45\"></td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"45\">Use this report to validate the benefit amounts that were calculated during payroll processing.</td>\n</tr>\n<tr sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"46\">\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"46\">Worker payment register</td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"46\">To comply with auditing best practices, use this report every pay period to validate data and sign off on pay runs.</td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"46\"></td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"46\"></td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"46\"></td>\n</tr>\n<tr sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"47\">\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"47\">Tax register</td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"47\">Use this report to validate the tax amounts that were calculated during payroll processing.</td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"47\">Use this report to validate the tax amounts that were calculated during payroll processing.</td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"47\">Use this report to validate the tax amounts that were calculated during payroll processing.</td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"47\">Use this report to validate the tax amounts that were calculated during payroll processing.</td>\n</tr>\n<tr sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"48\">\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"48\">State quarterly wage and tax preparation</td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"48\"></td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"48\">Use the information on this report when you prepare the quarterly wage and tax forms for state unemployment taxes.</td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"48\"></td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"48\"></td>\n</tr>\n<tr sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"49\">\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"49\">Form 941 preparation</td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"49\"></td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"49\">Use the information in this form when you prepare the quarterly report of payroll taxes for the Internal Revenue Service (IRS).</td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"49\"></td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"49\"></td>\n</tr>\n<tr sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"50\">\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"50\">Form 940 preparation</td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"50\"></td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"50\"></td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"50\">Use the information on this report when you prepare the annual federal unemployment tax (FUTA) return.</td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"50\"></td>\n</tr>\n<tr sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"51\">\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"51\">Form W-2 reconciliation</td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"51\"></td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"51\"></td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"51\">Use this report to balance Form W-2s and run validation before you issue Form W-2s to workers.</td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"51\">Use this report to balance Form W-2s and run validation before you issue Form W-2s to workers.</td>\n</tr>\n<tr sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"52\">\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"52\">Form W-2</td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"52\"></td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"52\"></td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"52\">Use this report to create Form W-2s that you can issue to workers.</td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"52\">Use this report to create Form W-2s that you can issue to workers.</td>\n</tr>\n<tr sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"53\">\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"53\">Electronic Form W-2</td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"53\"></td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"53\"></td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"53\">Use this report to file Form W-2s with the Social Security Administration.</td>\n<td sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"53\"></td>\n</tr>\n</tbody>\n</table>\n[!include[footer-include](../../../../includes/footer-banner.md)]","type":"Conceptual","source":{"$type":"Microsoft.DocAsCode.DataContracts.Common.SourceDetail, Microsoft.DocAsCode.DataContracts.Common","remote":{"$type":"Microsoft.DocAsCode.Common.Git.GitDetail, Microsoft.DocAsCode.Common","path":"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md","branch":"master","repo":"https://github.com/togoAIO/V0_DOKUD365.git"},"startLine":0,"endLine":0,"isExternal":false},"path":"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md","documentation":{"$type":"Microsoft.DocAsCode.DataContracts.Common.SourceDetail, Microsoft.DocAsCode.DataContracts.Common","remote":{"$type":"Microsoft.DocAsCode.Common.Git.GitDetail, Microsoft.DocAsCode.Common","path":"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md","branch":"master","repo":"https://github.com/togoAIO/V0_DOKUD365.git"},"startLine":0,"endLine":0,"isExternal":false},"_enableSearch":"true","_appFooter":"<span>Customized Footer</span>","_docfxVersion":"2.56.6.0","_appTitle":"WIKA Documentation","_systemKeys":{"$type":"System.String[], mscorlib","$values":["conceptual","type","source","path","documentation","title","rawTitle","wordCount"]},"rawTitle":"<h1 id=\"standard-payroll-reports\" sourcefile=\"ProcessDoku/02_SupportProcesses/02_01_Finance/hr/localizations/noam-usa-generate-payroll-reports.md\" sourcestartlinenumber=\"30\">Standard payroll reports</h1>","ms.custom":220994,"title":"Standard payroll reports","ms.dyn365.ops.version":"Version 1611","ms.search.region":"USA","ms.assetid":"92b0da78-1c42-46f7-b1a2-334d75e625f3","author":"andreabichsel","description":"This topic describes the standard payroll reports that are provided to help you with payroll processing and government reporting.","ms.author":"panolte","audience":"Application User","ms.search.validFrom":"2016-11-30","ms.topic":"article","ms.date":"06/20/2017","ms.technology":null,"ms.prod":null,"ms.reviewer":"anbichse"}�   �C  {"$type":"System.Collections.Generic.Dictionary`2[[System.String, mscorlib],[System.Object, mscorlib]], mscorlib","IsUserDefinedTitle":true,"XrefSpec":null}	   �C   